--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   17:11:02 10/23/2015
-- Design Name:   
-- Module Name:   C:/Experiments/mu2e/Readout_Controller/Controller_FPGA1/Controller_FPGA1_tb.vhd
-- Project Name:  Controller_FPGA1
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: ControllerFPGA_1
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use work.Project_defs.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

USE ieee.numeric_std.ALL;
library UNISIM;  

use UNISIM.Vcomponents.all;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;

ENTITY Controller_FPGA1_tb IS
END Controller_FPGA1_tb;

ARCHITECTURE behavior OF Controller_FPGA1_tb IS 

-- Component Declaration for the Unit Under Test (UUT)

 COMPONENT ControllerFPGA_1
 PORT
	(-- 159.3 MHz VXO clock, 50MHz Phy clock
	VXO_P,VXO_N,ClkB_P,ClkB_N,Clk50MHz,BnchClk : in std_logic;
-- 156.25 MHz GTP Reference clock, Gigabit data lines
	GTPClk_P,GTPClk_N,GTPRx_P,GTPRx_N : in std_logic_vector(1 downto 0);
	GTPTx_P,GTPTx_N : out std_logic_vector(1 downto 0);
-- Optical transcever slow control lines
	TDisA,TDisB : buffer std_logic;
--	SCLA,SDAA,SCLB,SDAB : inout std_logic;
	SD_A,SD_B : in std_logic;
-- microcontroller strobes
	CpldRst, CpldCS, uCRd, uCWr, EthCS : in std_logic;
-- microcontroller data, address buses
	uCA : in std_logic_vector(11 downto 0);
	uCD : inout std_logic_vector(15 downto 0);
-- Geographic address pins
	GA : in std_logic_vector(1 downto 0);
-- Serial inter-chip link clock, framing lines
	LINKClk_P,LINKClk_N,LinkFR_P,LinkFR_N  : in std_logic_vector(2 downto 0);
-- Serial inter-chip link Data lines
	LinkSDat_P,LinkSDat_N : in std_logic_vector(5 downto 0);
-- FM Transmitters for uBunch and Triggers
	HeartBeatFM,TrigFM,uBunchLED,TrigLED : buffer std_logic;
-- Pll control lines
	PllSClk,PllSDat,PllLd,PllPDn : buffer std_logic;
	PllStat : in std_logic;
-- Serial control lines for the RJ-45 LEDs
	LEDSClk,LEDSDat : out std_logic_vector(2 downto 0);
	LEDLd : out std_logic_vector(5 downto 0);
	LEDRst : buffer std_logic;
-- Orange Tree Ethernet daughter card lines
	DQ : inout std_logic_vector(15 downto 0);
	ZEthA : buffer std_logic_vector(8 downto 0);
	ZEthCS,ZEthWE,ZEthClk : buffer std_logic;
	ZEthBE : buffer std_logic_vector(1 downto 0);
	ZEthEOF : in std_logic_vector(1 downto 0);
	ZEthLen : in std_logic;
-- Back panel LEMOs
	GPO : buffer std_logic_vector(1 downto 0);
	GPI,NimTrig : in std_logic;
-- Debug port
	Debug : buffer std_logic_vector(10 downto 1));
	
 END COMPONENT;

signal VXO_P,VXO_N,ClkB_P,ClkB_N,Clk50MHz,BnchClk : std_logic;
signal GTPClk_P,GTPClk_N,GTPRx_P,GTPRx_N : std_logic_vector(1 downto 0);
signal GTPTx_P,GTPTx_N : std_logic_vector(1 downto 0);
signal TDisA,TDisB : std_logic;
signal SD_A,SD_B : std_logic;
signal CpldRst, CpldCS, uCRd, uCWr, EthCS : std_logic;
signal uCA : std_logic_vector(11 downto 0);
signal uCD : std_logic_vector(15 downto 0);
signal GA : std_logic_vector(1 downto 0);
signal LINKClk_P,LINKClk_N,LinkFR_P,LinkFR_N  : std_logic_vector(2 downto 0);
signal LinkSDat_P,LinkSDat_N : std_logic_vector(5 downto 0);
signal HeartBeatFM,TrigFM,uBunchLED,TrigLED : std_logic;
signal PllSClk,PllSDat,PllLd,PllPDn : std_logic;
signal PllStat : std_logic;
signal LEDSClk,LEDSDat : std_logic_vector(2 downto 0);
signal LEDLd : std_logic_vector(5 downto 0);
signal LEDRst : std_logic;
signal DQ : std_logic_vector(15 downto 0);
signal ZEthA : std_logic_vector(8 downto 0);
signal ZEthCS,ZEthWE,ZEthClk : std_logic;
signal ZEthBE : std_logic_vector(1 downto 0);
signal ZEthEOF : std_logic_vector(1 downto 0);
signal ZEthLen : std_logic;
signal GPO : std_logic_vector(1 downto 0);
signal GPI,NimTrig : std_logic;
signal Debug : std_logic_vector(10 downto 1);

-- Clock period definitions
constant ClkB_P_period : time := 6.25 ns; -- DG: NEW BOARD!!! 160MHz clock!!!
constant Clk53Mhz_Period : time := 18.83 ns;
constant DCO_period : time := 4 ns;
constant Clk50Mhz_Period : time := 20 ns;
constant Clk160Mhz_Period : time := 6.25 ns;
constant GTPRefClk_Period : time := 6.4 ns;
Constant GTP_Size : Integer := 48;

Type LEDTx_Array is Array(0 to GTP_Size - 1) of std_logic_vector(15 downto 0);
Constant TxVal : LEDTx_Array := (x"0000",x"0020",x"2345",x"3456",
                                 x"9210",x"0000",x"0000",x"0000",
											x"9122",x"9344",x"9566",x"9788",
                                 x"ABCC",x"ADEE",x"9F00",x"8003",
											x"1DED",x"8004",x"3AA9",x"8787",
											x"1122",x"3344",x"5566",x"7788",
                                 x"09AA",x"0BCC",x"3DEE",x"FF00",
											x"1DED",x"8004",x"3AA9",x"8787",
											x"1122",x"3344",x"5566",x"7788",
                                 x"09AA",x"3DEE",x"FF00",x"8004",
											x"1DED",x"2BCB",x"3AA9",x"8787",
                                 x"6565",x"4343",x"2121",x"8004");

Constant LinkDat0_Size : Integer := 221;
Type LinkDat0_Array is Array(0 to LinkDat0_Size - 1) of std_logic_vector(15 downto 0);
Constant LinkDat0 : LinkDat0_Array := 
(X"0004",X"0004",X"0000",X"0001",X"0100",X"0004",X"0000",X"0002",X"0100",
X"0004",X"0000",X"0003",X"0100",X"0004",X"0000",X"0004",X"0100",
X"0004",X"0000",X"0005",X"0100",X"0004",X"0000",X"0006",X"0100",
X"0004",X"0000",X"0007",X"0100",X"0004",X"0000",X"0008",X"0100",
X"0004",X"0000",X"0009",X"0100",X"0004",X"0000",X"000A",X"0100",
X"0004",X"0000",X"000B",X"0100",X"0004",X"0000",X"000C",X"0100",
X"0004",X"0000",X"000D",X"0100",X"0004",X"0000",X"000E",X"0100",
X"0004",X"0000",X"000F",X"0100",X"0004",X"0000",X"0010",X"0100",
X"0004",X"0000",X"0011",X"0100",X"0004",X"0000",X"0012",X"0100",
X"0004",X"0000",X"0013",X"0100",X"0004",X"0000",X"0014",X"0100",
X"0004",X"0000",X"0015",X"0100",X"0004",X"0000",X"0016",X"0100",
X"0004",X"0000",X"0017",X"0100",X"0004",X"0000",X"0018",X"0100",
X"0004",X"0000",X"0019",X"0100",X"0004",X"0000",X"001A",X"0100",
X"0004",X"0000",X"001B",X"0100",X"0004",X"0000",X"001C",X"0100",
X"0004",X"0000",X"001D",X"0100",X"0004",X"0000",X"001E",X"0100",
X"0004",X"0000",X"001F",X"0100",X"0004",X"0000",X"0020",X"0100",
X"0004",X"0000",X"0021",X"0100",X"0004",X"0000",X"0022",X"0100",
X"0004",X"0000",X"0023",X"0100",X"0004",X"0000",X"0024",X"0100",
X"0004",X"0000",X"0025",X"0100",X"0004",X"0000",X"0026",X"0100",
X"0004",X"0000",X"0027",X"0100",X"0004",X"0000",X"0028",X"0100",
X"000E",X"0000",X"0029",X"0100",X"0018",X"4005",X"0007",X"002C",
X"0006",X"0FE2",X"0FE7",X"0FF4",X"0FF8",X"0FF7",X"0004",X"0000",
X"002A",X"0100",X"0004",X"0000",X"002B",X"0100",X"0004",X"0000",
X"002C",X"0100",X"0004",X"0000",X"002D",X"0100",X"000E",X"0000",
X"002E",X"0100",X"0018",X"4012",X"0FF9",X"0019",X"0027",X"0FF7",
X"0FE0",X"0FEA",X"0FF8",X"0FF7",X"0004",X"0000",X"002F",X"0100",
X"0004",X"0000",X"0030",X"0100",X"0004",X"0000",X"0031",X"0100",
X"0004",X"0000",X"0000",X"0100");

--Constant LinkDat0_Size : Integer := 5586;
--Type LinkDat0_Array is Array(0 to LinkDat0_Size - 1) of std_logic_vector(15 downto 0);
--Constant LinkDat0 : LinkDat0_Array := 
--(X"01E8",X"01E8",X"FF00",X"0060",X"0042",X"0000",X"FFFF",X"03E8",X"0000",
--X"FF01",X"FF00",X"0004",X"03E8",X"0008",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0033",X"03E8",X"000A",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"00E0",X"0030",X"03E8",X"0005",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0016",X"03E8",X"0003",X"00BB",X"0164",X"06DB",
--X"0004",X"03E8",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"000A",X"03E8",X"0006",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"0060",X"0059",X"0001",X"FFFF",
--X"03E8",X"0000",X"FF01",X"FF00",X"0057",X"03E8",X"0003",X"00BB",
--X"0164",X"06DB",X"0049",X"03E8",X"0004",X"00BB",X"0164",X"06DB",
--X"0F1B",X"007C",X"03E8",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0068",X"03E8",X"0003",X"00BB",X"0164",X"06DB",X"0063",
--X"03E8",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"012A",X"006A",X"03E8",X"0003",X"00BB",X"0164",
--X"06DB",X"0069",X"03E8",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0078",X"03E8",
--X"0003",X"00BB",X"0164",X"06DB",X"0052",X"03E8",X"0004",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0042",X"03E8",X"0007",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0060",X"0028",X"0002",
--X"FFFF",X"03E8",X"0000",X"FF01",X"FF00",X"0099",X"03E8",X"0004",
--X"00BB",X"0164",X"06DB",X"0F1B",X"00A9",X"03E8",X"0005",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"008A",X"03E8",X"0008",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0098",
--X"03E8",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"0065",X"0003",
--X"FFFF",X"03E8",X"0000",X"FF01",X"FF00",X"00E9",X"03E8",X"0003",
--X"00BB",X"0164",X"06DB",X"00E1",X"03E8",X"0008",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"00E9",X"03E8",
--X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00E6",X"03E8",X"0005",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"00EE",X"03E8",X"0004",X"00BB",X"0164",X"06DB",
--X"0F1B",X"00F1",X"03E8",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
--X"00F1",X"03E8",X"0003",X"00BB",X"0164",X"06DB",X"00E9",X"03E8",
--X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00E0",X"00CD",X"03E8",X"0008",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"00E0",X"03E8",
--X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"0060",X"0022",X"0004",X"FFFF",X"03E8",X"0000",
--X"FF01",X"FF00",X"0033",X"03E8",X"0004",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0012",X"03E8",X"0003",X"00BB",X"0164",X"06DB",X"0022",
--X"03E8",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"012A",X"00E0",X"0060",X"0036",X"0005",X"FFFF",
--X"03E8",X"0000",X"FF01",X"FF00",X"005D",X"03E8",X"0003",X"00BB",
--X"0164",X"06DB",X"006C",X"03E8",X"0008",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0076",X"03E8",X"000A",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"00E0",X"0060",X"03E8",X"0007",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"007F",X"03E8",X"0003",X"00BB",
--X"0164",X"06DB",X"0060",X"004D",X"0006",X"FFFF",X"03E8",X"0000",
--X"FF01",X"FF00",X"0099",X"03E8",X"0003",X"00BB",X"0164",X"06DB",
--X"00AA",X"03E8",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0099",X"03E8",X"0008",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"00A0",X"03E8",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"00B6",X"03E8",X"0006",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"0082",X"03E8",X"0005",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0087",X"03E8",X"0008",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0060",
--X"0019",X"0007",X"FFFF",X"03E8",X"0000",X"FF01",X"FF00",X"00DF",
--X"03E8",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"00E5",X"03E8",X"0003",X"00BB",X"0164",X"06DB",
--X"01F7",X"FF00",X"0060",X"0027",X"0000",X"FFFF",X"03F2",X"0001",
--X"FF01",X"FF00",X"0006",X"03F2",X"0006",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"002A",X"03F2",X"0005",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0004",X"03F2",X"0005",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0002",X"03F2",X"0003",X"00BB",X"0164",
--X"06DB",X"0060",X"006A",X"0001",X"FFFF",X"03F2",X"0001",X"FF01",
--X"FF00",X"0042",X"03F2",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"006B",X"03F2",X"0009",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"004F",
--X"03F2",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"007B",X"03F2",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"0055",X"03F2",X"0006",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0059",X"03F2",X"0006",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0060",X"03F2",
--X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0069",X"03F2",X"0006",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"004F",X"03F2",
--X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0071",X"03F2",
--X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00E0",X"0060",X"004D",X"0002",X"FFFF",X"03F2",
--X"0001",X"FF01",X"FF00",X"008D",X"03F2",X"0007",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"00A1",X"03F2",X"0003",
--X"00BB",X"0164",X"06DB",X"00B6",X"03F2",X"000A",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
--X"009E",X"03F2",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"00A7",X"03F2",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"00B7",X"03F2",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"00E0",X"008D",X"03F2",X"0008",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"0060",X"0008",X"0003",X"FFFF",X"03F2",X"0001",X"FF01",X"FF00",
--X"0060",X"000E",X"0004",X"FFFF",X"03F2",X"0001",X"FF01",X"FF00",
--X"0006",X"03F2",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"005B",
--X"0005",X"FFFF",X"03F2",X"0001",X"FF01",X"FF00",X"0075",X"03F2",
--X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"004C",X"03F2",X"0005",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0042",X"03F2",X"0007",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"006C",X"03F2",X"0007",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"007A",X"03F2",
--X"0003",X"00BB",X"0164",X"06DB",X"0049",X"03F2",X"0006",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"006A",X"03F2",X"0005",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"006C",X"03F2",X"0007",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"004B",
--X"03F2",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"0060",X"0053",X"0006",X"FFFF",X"03F2",X"0001",X"FF01",
--X"FF00",X"00A4",X"03F2",X"0003",X"00BB",X"0164",X"06DB",X"0099",
--X"03F2",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"012A",X"00A5",X"03F2",X"0004",X"00BB",X"0164",
--X"06DB",X"0F1B",X"009F",X"03F2",X"0006",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"0083",X"03F2",X"0004",X"00BB",X"0164",
--X"06DB",X"0F1B",X"009B",X"03F2",X"0005",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"00A8",X"03F2",X"0003",X"00BB",X"0164",X"06DB",
--X"008C",X"03F2",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"008D",X"03F2",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"0060",X"0053",X"0007",X"FFFF",
--X"03F2",X"0001",X"FF01",X"FF00",X"00D4",X"03F2",X"0003",X"00BB",
--X"0164",X"06DB",X"00C5",X"03F2",X"0008",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"00FB",X"03F2",X"0008",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"00C7",X"03F2",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"00F7",X"03F2",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"00FD",X"03F2",X"0004",
--X"00BB",X"0164",X"06DB",X"0F1B",X"00F5",X"03F2",X"0008",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"00E7",
--X"03F2",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"01AA",
--X"FF00",X"0060",X"0008",X"0000",X"FFFF",X"03FC",X"0002",X"FF01",
--X"FF00",X"0060",X"0060",X"0001",X"FFFF",X"03FC",X"0002",X"FF01",
--X"FF00",X"005A",X"03FC",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"004E",X"03FC",X"0006",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0054",X"03FC",X"0008",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"0073",X"03FC",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"0040",X"03FC",X"0009",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
--X"007C",X"03FC",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0069",
--X"03FC",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"007B",X"03FC",
--X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"004D",X"03FC",X"0004",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0060",X"001B",X"0002",X"FFFF",X"03FC",X"0002",X"FF01",
--X"FF00",X"008C",X"03FC",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"00A6",X"03FC",
--X"0003",X"00BB",X"0164",X"06DB",X"0060",X"0024",X"0003",X"FFFF",
--X"03FC",X"0002",X"FF01",X"FF00",X"00D0",X"03FC",X"0004",X"00BB",
--X"0164",X"06DB",X"0F1B",X"00D3",X"03FC",X"0006",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"00C5",X"03FC",X"0009",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
--X"0060",X"0038",X"0004",X"FFFF",X"03FC",X"0002",X"FF01",X"FF00",
--X"0008",X"03FC",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0004",X"03FC",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"0019",X"03FC",X"0004",X"00BB",
--X"0164",X"06DB",X"0F1B",X"002D",X"03FC",X"0008",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"003A",X"03FC",
--X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"0060",X"0042",X"0005",X"FFFF",X"03FC",X"0002",X"FF01",X"FF00",
--X"0043",X"03FC",X"0003",X"00BB",X"0164",X"06DB",X"005E",X"03FC",
--X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"0045",X"03FC",X"0009",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0040",X"03FC",
--X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0056",X"03FC",
--X"0003",X"00BB",X"0164",X"06DB",X"0071",X"03FC",X"0003",X"00BB",
--X"0164",X"06DB",X"0061",X"03FC",X"0005",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0060",X"0038",X"0006",X"FFFF",X"03FC",X"0002",
--X"FF01",X"FF00",X"0091",X"03FC",X"0009",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00AF",X"03FC",
--X"0003",X"00BB",X"0164",X"06DB",X"0087",X"03FC",X"000A",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
--X"00E0",X"00AC",X"03FC",X"0003",X"00BB",X"0164",X"06DB",X"009A",
--X"03FC",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"0060",X"004F",X"0007",X"FFFF",X"03FC",X"0002",
--X"FF01",X"FF00",X"00F0",X"03FC",X"0006",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"00FC",X"03FC",X"0008",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"00F7",X"03FC",
--X"0003",X"00BB",X"0164",X"06DB",X"00D6",X"03FC",X"0005",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"00C2",X"03FC",X"0006",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"00F8",X"03FC",X"0006",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"00D9",X"03FC",
--X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"00D9",
--X"03FC",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01D1",X"FF00",X"0060",X"0008",X"0000",X"FFFF",X"0406",
--X"0003",X"FF01",X"FF00",X"0060",X"0066",X"0001",X"FFFF",X"0406",
--X"0003",X"FF01",X"FF00",X"0062",X"0406",X"0007",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0044",X"0406",X"0006",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0069",X"0406",
--X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"0046",X"0406",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"0055",X"0406",X"0009",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"007D",
--X"0406",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"006F",X"0406",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"007E",X"0406",X"0005",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0044",X"0406",X"0009",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"0060",X"000E",X"0002",X"FFFF",X"0406",X"0003",X"FF01",
--X"FF00",X"009F",X"0406",X"0003",X"00BB",X"0164",X"06DB",X"0060",
--X"0032",X"0003",X"FFFF",X"0406",X"0003",X"FF01",X"FF00",X"00FA",
--X"0406",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"00F0",X"0406",X"0005",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"00DF",X"0406",X"0007",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"00D0",X"0406",X"000A",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
--X"00E0",X"0060",X"003E",X"0004",X"FFFF",X"0406",X"0003",X"FF01",
--X"FF00",X"0035",X"0406",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"003C",X"0406",
--X"0003",X"00BB",X"0164",X"06DB",X"001D",X"0406",X"000A",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
--X"00E0",X"0009",X"0406",X"0003",X"00BB",X"0164",X"06DB",X"0032",
--X"0406",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"0024",X"0406",X"0003",X"00BB",X"0164",X"06DB",X"0060",
--X"004B",X"0005",X"FFFF",X"0406",X"0003",X"FF01",X"FF00",X"007F",
--X"0406",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"0066",X"0406",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"0062",X"0406",X"000A",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
--X"00E0",X"0072",X"0406",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"006E",X"0406",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"004C",X"0406",X"000A",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"00E0",X"0060",X"0044",X"0006",X"FFFF",X"0406",X"0003",
--X"FF01",X"FF00",X"009A",X"0406",X"0005",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"00AF",X"0406",X"0006",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"009C",X"0406",X"0008",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0083",X"0406",
--X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"00B2",X"0406",X"0003",
--X"00BB",X"0164",X"06DB",X"00B1",X"0406",X"0003",X"00BB",X"0164",
--X"06DB",X"009A",X"0406",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0060",X"0054",
--X"0007",X"FFFF",X"0406",X"0003",X"FF01",X"FF00",X"00FC",X"0406",
--X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"00F3",X"0406",
--X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"00E1",X"0406",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"00C4",X"0406",X"0004",X"00BB",
--X"0164",X"06DB",X"0F1B",X"00E4",X"0406",X"000A",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
--X"00E9",X"0406",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"00D0",X"0406",X"0004",X"00BB",X"0164",
--X"06DB",X"0F1B",X"00CC",X"0406",X"0005",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"023B",X"FF00",X"0060",X"003B",X"0000",X"FFFF",
--X"0410",X"0004",X"FF01",X"FF00",X"0035",X"0410",X"0009",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
--X"0013",X"0410",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"0023",X"0410",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0034",X"0410",
--X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0000",X"0410",
--X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0060",
--X"0063",X"0001",X"FFFF",X"0410",X"0004",X"FF01",X"FF00",X"0077",
--X"0410",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0046",X"0410",
--X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0074",
--X"0410",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"004F",X"0410",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0079",X"0410",X"0003",
--X"00BB",X"0164",X"06DB",X"0073",X"0410",X"0006",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"0047",X"0410",X"000A",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
--X"00E0",X"004D",X"0410",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
--X"006D",X"0410",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"0073",X"0410",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"0060",X"0025",X"0002",X"FFFF",X"0410",X"0004",
--X"FF01",X"FF00",X"00B1",X"0410",X"0008",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"00A3",X"0410",X"0003",
--X"00BB",X"0164",X"06DB",X"00B7",X"0410",X"0009",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0060",
--X"0064",X"0003",X"FFFF",X"0410",X"0004",X"FF01",X"FF00",X"00D2",
--X"0410",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"00F6",X"0410",X"0008",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"00DA",X"0410",X"0007",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"00EC",
--X"0410",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"00CA",X"0410",X"0003",X"00BB",X"0164",X"06DB",X"00D9",X"0410",
--X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"00DE",X"0410",X"0009",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"00FB",X"0410",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"00E1",X"0410",X"0006",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"00C1",X"0410",X"0004",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0060",X"0054",X"0004",X"FFFF",X"0410",
--X"0004",X"FF01",X"FF00",X"0010",X"0410",X"000A",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
--X"000C",X"0410",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"00E0",X"003B",X"0410",X"0004",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0021",X"0410",X"0007",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"003F",X"0410",
--X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00E0",X"0030",X"0410",X"0005",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0029",X"0410",X"0009",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0060",
--X"001D",X"0005",X"FFFF",X"0410",X"0004",X"FF01",X"FF00",X"006C",
--X"0410",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"006F",X"0410",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"0060",X"0072",X"0006",X"FFFF",
--X"0410",X"0004",X"FF01",X"FF00",X"0082",X"0410",X"0008",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0092",
--X"0410",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"008E",X"0410",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"00BE",X"0410",X"0006",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"009B",X"0410",X"000A",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
--X"0092",X"0410",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0087",X"0410",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"00E0",X"00BB",X"0410",X"0005",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"00BC",X"0410",X"0009",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"008D",X"0410",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0060",X"002F",
--X"0007",X"FFFF",X"0410",X"0004",X"FF01",X"FF00",X"00EB",X"0410",
--X"0003",X"00BB",X"0164",X"06DB",X"00E8",X"0410",X"0005",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"00D7",X"0410",X"0003",X"00BB",
--X"0164",X"06DB",X"00C1",X"0410",X"0008",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"00EB",X"0410",X"0005",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"018C",X"FF00",X"0060",
--X"0022",X"0000",X"FFFF",X"041A",X"0005",X"FF01",X"FF00",X"0006",
--X"041A",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"012A",X"001F",X"041A",X"0003",X"00BB",X"0164",
--X"06DB",X"0018",X"041A",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0060",X"0008",X"0001",X"FFFF",X"041A",X"0005",X"FF01",
--X"FF00",X"0060",X"0047",X"0002",X"FFFF",X"041A",X"0005",X"FF01",
--X"FF00",X"00B8",X"041A",X"0003",X"00BB",X"0164",X"06DB",X"00AF",
--X"041A",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"012A",X"008C",X"041A",X"0004",X"00BB",X"0164",
--X"06DB",X"0F1B",X"00B0",X"041A",X"0006",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"008C",X"041A",X"0009",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0097",
--X"041A",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"00B7",
--X"041A",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"0060",X"003C",X"0003",X"FFFF",X"041A",X"0005",X"FF01",X"FF00",
--X"00D1",X"041A",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"00D9",X"041A",X"0005",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"00E5",X"041A",X"0007",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"00D3",X"041A",X"0009",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"00E6",X"041A",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"0060",X"001F",X"0004",X"FFFF",
--X"041A",X"0005",X"FF01",X"FF00",X"0004",X"041A",X"0009",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
--X"0035",X"041A",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"0060",X"0040",X"0005",X"FFFF",X"041A",
--X"0005",X"FF01",X"FF00",X"0049",X"041A",X"0006",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"0075",X"041A",X"000A",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
--X"00E0",X"0047",X"041A",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"0054",X"041A",X"000A",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"00E0",X"005E",X"041A",X"0006",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"0060",X"0040",X"0006",X"FFFF",X"041A",
--X"0005",X"FF01",X"FF00",X"00A9",X"041A",X"0006",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"00A5",X"041A",X"0009",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
--X"0092",X"041A",X"0003",X"00BB",X"0164",X"06DB",X"00B6",X"041A",
--X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"00B3",X"041A",
--X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"00B5",X"041A",
--X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00E0",X"0060",X"003E",X"0007",X"FFFF",X"041A",
--X"0005",X"FF01",X"FF00",X"00CA",X"041A",X"0004",X"00BB",X"0164",
--X"06DB",X"0F1B",X"00F9",X"041A",X"0005",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"00E1",X"041A",X"0009",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00F1",X"041A",
--X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"00C7",X"041A",X"000A",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"00E0",X"00C4",X"041A",X"0004",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0220",X"FF00",X"0060",X"0008",X"0000",X"FFFF",X"0424",
--X"0006",X"FF01",X"FF00",X"0060",X"003A",X"0001",X"FFFF",X"0424",
--X"0006",X"FF01",X"FF00",X"0058",X"0424",X"0007",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0059",X"0424",X"0009",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"007A",X"0424",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0077",X"0424",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"0063",X"0424",X"0007",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0060",X"0039",X"0002",
--X"FFFF",X"0424",X"0006",X"FF01",X"FF00",X"0088",X"0424",X"0009",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"0091",X"0424",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"009A",X"0424",
--X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00E0",X"0093",X"0424",X"0008",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0060",X"005E",
--X"0003",X"FFFF",X"0424",X"0006",X"FF01",X"FF00",X"00E3",X"0424",
--X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"00FC",X"0424",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"00E0",X"00D7",X"0424",X"0006",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"00E3",X"0424",
--X"0003",X"00BB",X"0164",X"06DB",X"00C8",X"0424",X"0008",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"00CE",
--X"0424",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"00E5",X"0424",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"00F3",X"0424",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
--X"00E1",X"0424",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"0060",X"003C",X"0004",X"FFFF",
--X"0424",X"0006",X"FF01",X"FF00",X"0022",X"0424",X"0004",X"00BB",
--X"0164",X"06DB",X"0F1B",X"000A",X"0424",X"0007",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0014",X"0424",X"0004",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0033",X"0424",X"0005",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"000C",X"0424",X"0007",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"000E",X"0424",
--X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"0060",X"004C",X"0005",X"FFFF",X"0424",X"0006",X"FF01",X"FF00",
--X"0063",X"0424",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"004E",
--X"0424",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0049",X"0424",
--X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"0055",X"0424",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"0074",X"0424",X"0008",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0053",X"0424",
--X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"004F",
--X"0424",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"012A",X"00E0",X"0060",X"005A",X"0006",X"FFFF",
--X"0424",X"0006",X"FF01",X"FF00",X"008B",X"0424",X"0003",X"00BB",
--X"0164",X"06DB",X"009A",X"0424",X"0006",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"00B2",X"0424",X"0006",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"008C",X"0424",X"0005",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"00A4",X"0424",X"0007",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"00A2",X"0424",
--X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"00B0",X"0424",
--X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"00B4",
--X"0424",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"00A1",X"0424",X"0003",X"00BB",X"0164",X"06DB",
--X"00A5",X"0424",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"0063",
--X"0007",X"FFFF",X"0424",X"0006",X"FF01",X"FF00",X"00FE",X"0424",
--X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"00C3",
--X"0424",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"00E5",X"0424",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"00C7",X"0424",X"0004",X"00BB",X"0164",X"06DB",
--X"0F1B",X"00D6",X"0424",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"00E3",X"0424",X"000A",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
--X"00D9",X"0424",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"00CE",X"0424",X"0007",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"00C1",X"0424",X"0009",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"01D9",X"FF00",X"0060",X"0032",X"0000",X"FFFF",X"042E",
--X"0007",X"FF01",X"FF00",X"0027",X"042E",X"0004",X"00BB",X"0164",
--X"06DB",X"0F1B",X"003E",X"042E",X"000A",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0028",
--X"042E",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"0009",X"042E",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0060",X"003E",X"0001",
--X"FFFF",X"042E",X"0007",X"FF01",X"FF00",X"004A",X"042E",X"0007",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0070",
--X"042E",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"005F",X"042E",X"0004",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0071",X"042E",X"0003",X"00BB",X"0164",X"06DB",X"0050",
--X"042E",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"005B",X"042E",
--X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00E0",X"0060",X"000E",X"0002",X"FFFF",X"042E",
--X"0007",X"FF01",X"FF00",X"00A1",X"042E",X"0003",X"00BB",X"0164",
--X"06DB",X"0060",X"003E",X"0003",X"FFFF",X"042E",X"0007",X"FF01",
--X"FF00",X"00D6",X"042E",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"00FC",X"042E",
--X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00D8",X"042E",X"0003",X"00BB",X"0164",X"06DB",
--X"00C7",X"042E",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"00E6",
--X"042E",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"00E6",X"042E",
--X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0060",
--X"003E",X"0004",X"FFFF",X"042E",X"0007",X"FF01",X"FF00",X"0002",
--X"042E",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"0036",X"042E",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"002C",X"042E",X"0005",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0004",X"042E",X"0004",X"00BB",X"0164",X"06DB",
--X"0F1B",X"001C",X"042E",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0035",X"042E",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"0060",X"002C",X"0005",
--X"FFFF",X"042E",X"0007",X"FF01",X"FF00",X"004D",X"042E",X"0009",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"007E",X"042E",X"0003",X"00BB",X"0164",X"06DB",X"0064",
--X"042E",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"0050",X"042E",X"0004",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0060",X"0049",X"0006",X"FFFF",X"042E",X"0007",X"FF01",
--X"FF00",X"00B4",X"042E",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"00AF",X"042E",X"000A",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
--X"00B3",X"042E",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"00E0",X"00AD",X"042E",X"0007",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0084",
--X"042E",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"009E",X"042E",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"0060",X"0068",X"0007",X"FFFF",X"042E",X"0007",
--X"FF01",X"FF00",X"00D0",X"042E",X"0006",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"00CC",X"042E",X"0007",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"00DB",X"042E",X"0008",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"00C0",X"042E",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"00E6",X"042E",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"00DD",X"042E",X"0005",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"00FC",X"042E",X"0008",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"00DC",
--X"042E",X"0003",X"00BB",X"0164",X"06DB",X"00DC",X"042E",X"0007",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"00CE",
--X"042E",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"0178",X"FF00",X"0060",X"003A",X"0000",X"FFFF",
--X"0438",X"0008",X"FF01",X"FF00",X"0009",X"0438",X"0006",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"000B",X"0438",X"0005",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"003D",X"0438",X"000A",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"00E0",X"0033",X"0438",X"0008",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0014",X"0438",X"0006",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0060",X"0022",
--X"0001",X"FFFF",X"0438",X"0008",X"FF01",X"FF00",X"005B",X"0438",
--X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00E0",X"0063",X"0438",X"000A",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
--X"0060",X"0065",X"0002",X"FFFF",X"0438",X"0008",X"FF01",X"FF00",
--X"0093",X"0438",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"00B2",X"0438",X"0007",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"00B3",X"0438",X"0006",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0080",X"0438",
--X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"00B2",X"0438",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"00BD",X"0438",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"0098",X"0438",X"0007",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"00A5",X"0438",
--X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"008E",X"0438",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0060",X"0030",X"0003",
--X"FFFF",X"0438",X"0008",X"FF01",X"FF00",X"00EB",X"0438",X"0003",
--X"00BB",X"0164",X"06DB",X"00F8",X"0438",X"0009",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E4",
--X"0438",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"00CE",X"0438",X"0008",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0060",X"0013",X"0004",
--X"FFFF",X"0438",X"0008",X"FF01",X"FF00",X"002C",X"0438",X"0008",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"0060",X"0013",X"0005",X"FFFF",X"0438",X"0008",X"FF01",X"FF00",
--X"0049",X"0438",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"0060",X"0008",X"0006",X"FFFF",X"0438",
--X"0008",X"FF01",X"FF00",X"0060",X"0057",X"0007",X"FFFF",X"0438",
--X"0008",X"FF01",X"FF00",X"00C5",X"0438",X"000A",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
--X"00E6",X"0438",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"00F6",X"0438",X"0007",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"00FC",X"0438",X"0009",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
--X"00EA",X"0438",X"0003",X"00BB",X"0164",X"06DB",X"00C7",X"0438",
--X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"00E1",X"0438",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
--X"00CA",X"0438",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"0178",X"FF00",X"0060",X"0044",X"0000",X"FFFF",
--X"0442",X"0009",X"FF01",X"FF00",X"0037",X"0442",X"0007",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0035",X"0442",
--X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"0006",X"0442",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0029",X"0442",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0006",X"0442",X"0003",X"00BB",X"0164",X"06DB",X"001D",X"0442",
--X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0037",X"0442",
--X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"0060",X"000F",X"0001",X"FFFF",X"0442",X"0009",X"FF01",X"FF00",
--X"0050",X"0442",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0060",
--X"0015",X"0002",X"FFFF",X"0442",X"0009",X"FF01",X"FF00",X"0099",
--X"0442",X"0003",X"00BB",X"0164",X"06DB",X"00B9",X"0442",X"0004",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0060",X"005F",X"0003",X"FFFF",
--X"0442",X"0009",X"FF01",X"FF00",X"00C6",X"0442",X"0005",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"00C6",X"0442",X"000A",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
--X"00E0",X"00DA",X"0442",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"00CF",X"0442",
--X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"00CE",X"0442",
--X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00E9",X"0442",X"0003",X"00BB",X"0164",X"06DB",
--X"00CE",X"0442",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"00D1",X"0442",X"0006",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"00F5",X"0442",X"0003",
--X"00BB",X"0164",X"06DB",X"0060",X"0050",X"0004",X"FFFF",X"0442",
--X"0009",X"FF01",X"FF00",X"0038",X"0442",X"0004",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0037",X"0442",X"0007",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"000F",X"0442",X"0009",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
--X"000A",X"0442",X"0003",X"00BB",X"0164",X"06DB",X"0013",X"0442",
--X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00E0",X"000E",X"0442",X"0009",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0010",
--X"0442",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"012A",X"0060",X"0048",X"0005",X"FFFF",X"0442",
--X"0009",X"FF01",X"FF00",X"0077",X"0442",X"000A",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
--X"0058",X"0442",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"007B",X"0442",X"0003",X"00BB",
--X"0164",X"06DB",X"0053",X"0442",X"0005",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0064",X"0442",X"0009",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0046",X"0442",
--X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00E0",X"0060",X"0008",X"0006",X"FFFF",X"0442",
--X"0009",X"FF01",X"FF00",X"0060",X"000F",X"0007",X"FFFF",X"0442",
--X"0009",X"FF01",X"FF00",X"00DA",X"0442",X"0004",X"00BB",X"0164",
--X"06DB",X"0F1B",X"018E",X"FF00",X"0060",X"0050",X"0000",X"FFFF",
--X"044C",X"000A",X"FF01",X"FF00",X"002B",X"044C",X"0008",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0032",
--X"044C",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"001D",X"044C",X"0003",X"00BB",X"0164",X"06DB",
--X"001A",X"044C",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"0006",X"044C",X"0004",X"00BB",X"0164",
--X"06DB",X"0F1B",X"001B",X"044C",X"0003",X"00BB",X"0164",X"06DB",
--X"0028",X"044C",X"0003",X"00BB",X"0164",X"06DB",X"003B",X"044C",
--X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"002A",X"044C",
--X"0003",X"00BB",X"0164",X"06DB",X"0060",X"0015",X"0001",X"FFFF",
--X"044C",X"000A",X"FF01",X"FF00",X"0057",X"044C",X"0004",X"00BB",
--X"0164",X"06DB",X"0F1B",X"006A",X"044C",X"0003",X"00BB",X"0164",
--X"06DB",X"0060",X"003C",X"0002",X"FFFF",X"044C",X"000A",X"FF01",
--X"FF00",X"00B7",X"044C",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"00A3",X"044C",X"0009",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"0088",X"044C",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"00A8",X"044C",X"0003",
--X"00BB",X"0164",X"06DB",X"008E",X"044C",X"0007",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0060",X"0068",X"0003",
--X"FFFF",X"044C",X"000A",X"FF01",X"FF00",X"00C9",X"044C",X"0009",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"00F3",X"044C",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
--X"00F6",X"044C",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"00CD",X"044C",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"00DB",X"044C",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"00CC",X"044C",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"00C7",X"044C",X"0005",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"00E2",X"044C",X"0005",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"00EF",X"044C",X"000A",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"00E0",X"00F1",X"044C",X"0008",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0060",X"002B",X"0004",
--X"FFFF",X"044C",X"000A",X"FF01",X"FF00",X"0027",X"044C",X"0009",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"002D",X"044C",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"0032",X"044C",X"0008",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"0060",X"001A",X"0005",X"FFFF",X"044C",X"000A",X"FF01",X"FF00",
--X"0057",X"044C",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"0065",X"044C",X"0004",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0060",X"0008",X"0006",X"FFFF",X"044C",X"000A",
--X"FF01",X"FF00",X"0060",X"0036",X"0007",X"FFFF",X"044C",X"000A",
--X"FF01",X"FF00",X"00C6",X"044C",X"0004",X"00BB",X"0164",X"06DB",
--X"0F1B",X"00CC",X"044C",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"00C7",X"044C",
--X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00E0",X"00F0",X"044C",X"000A",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
--X"0239",X"FF00",X"0060",X"0019",X"0000",X"FFFF",X"0456",X"000B",
--X"FF01",X"FF00",X"0005",X"0456",X"0003",X"00BB",X"0164",X"06DB",
--X"0037",X"0456",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"0060",X"000E",X"0001",X"FFFF",X"0456",
--X"000B",X"FF01",X"FF00",X"007F",X"0456",X"0003",X"00BB",X"0164",
--X"06DB",X"0060",X"0064",X"0002",X"FFFF",X"0456",X"000B",X"FF01",
--X"FF00",X"0083",X"0456",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"012A",X"0087",X"0456",X"000A",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"00E0",X"00AA",X"0456",X"0007",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"00BD",X"0456",X"0008",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0085",
--X"0456",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0096",X"0456",
--X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"008B",X"0456",X"0003",X"00BB",X"0164",X"06DB",X"00BF",X"0456",
--X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00A2",X"0456",X"0008",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0060",X"0047",X"0003",
--X"FFFF",X"0456",X"000B",X"FF01",X"FF00",X"00E7",X"0456",X"0003",
--X"00BB",X"0164",X"06DB",X"00D6",X"0456",X"0008",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"00C4",X"0456",
--X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"00C6",X"0456",
--X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"00C6",X"0456",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"00C8",X"0456",X"0003",X"00BB",X"0164",
--X"06DB",X"00DD",X"0456",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"0060",X"004F",X"0004",X"FFFF",
--X"0456",X"000B",X"FF01",X"FF00",X"0025",X"0456",X"0007",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"000C",X"0456",
--X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"001E",X"0456",X"0004",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0002",X"0456",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"0032",X"0456",X"0007",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0004",X"0456",
--X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0028",X"0456",
--X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00E0",X"0060",X"003B",X"0005",X"FFFF",X"0456",
--X"000B",X"FF01",X"FF00",X"007A",X"0456",X"0007",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"005F",X"0456",X"000A",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"00E0",X"0077",X"0456",X"0003",X"00BB",X"0164",X"06DB",
--X"0050",X"0456",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"0064",X"0456",X"0008",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0060",X"0068",
--X"0006",X"FFFF",X"0456",X"000B",X"FF01",X"FF00",X"0092",X"0456",
--X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00E0",X"0083",X"0456",X"0008",X"00BB",X"0164",
--X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"00AE",X"0456",
--X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00B9",X"0456",X"0003",X"00BB",X"0164",X"06DB",
--X"0091",X"0456",X"0003",X"00BB",X"0164",X"06DB",X"0099",X"0456",
--X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"008B",X"0456",X"000A",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"00B0",
--X"0456",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C",X"01E3",X"00AA",X"0456",X"0009",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0060",X"0073",
--X"0007",X"FFFF",X"0456",X"000B",X"FF01",X"FF00",X"00E7",X"0456",
--X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"00C8",
--X"0456",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"00DC",X"0456",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
--X"0607",X"036C",X"01E3",X"012A",X"00C3",X"0456",X"0006",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"00FE",X"0456",X"0009",
--X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
--X"012A",X"00C1",X"0456",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
--X"0980",X"0607",X"036C",X"01E3",X"00EA",X"0456",X"0007",X"00BB",
--X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"00C5",X"0456",
--X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
--X"01E3",X"012A",X"00E8",X"0456",X"000A",X"00BB",X"0164",X"06DB",
--X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"00F5",
--X"0456",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
--X"036C");

Constant LinkDat1_Size : Integer := 5351;
Type LinkDat1_Array is Array(0 to LinkDat1_Size - 1) of std_logic_vector(15 downto 0);
Constant LinkDat1 : LinkDat1_Array := 
(X"01E8",X"01FD",X"FF00",X"0060",X"0042",X"0008",X"FFFF",X"03E8",X"0000",
X"FF01",X"FF00",X"020B",X"03E8",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"0231",X"03E8",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
X"0228",X"03E8",X"0003",X"00BB",X"0164",X"06DB",X"023F",X"03E8",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0201",X"03E8",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"021F",
X"03E8",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"020F",
X"03E8",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"0060",X"0048",X"0009",X"FFFF",
X"03E8",X"0000",X"FF01",X"FF00",X"026E",X"03E8",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"0261",X"03E8",X"0003",X"00BB",X"0164",X"06DB",X"0256",X"03E8",
X"0003",X"00BB",X"0164",X"06DB",X"0256",X"03E8",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0252",X"03E8",
X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"025D",X"03E8",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"024D",X"03E8",X"0007",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"0060",X"0020",X"000A",X"FFFF",
X"03E8",X"0000",X"FF01",X"FF00",X"02AD",X"03E8",X"0005",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"02A4",X"03E8",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0297",X"03E8",
X"0003",X"00BB",X"0164",X"06DB",X"0060",X"005A",X"000B",X"FFFF",
X"03E8",X"0000",X"FF01",X"FF00",X"02E7",X"03E8",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"02D6",X"03E8",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"02D7",X"03E8",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"02CD",X"03E8",X"0003",
X"00BB",X"0164",X"06DB",X"02D3",X"03E8",X"0005",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"02FE",X"03E8",X"0009",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"02FF",
X"03E8",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"02F5",X"03E8",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0060",X"002E",
X"000C",X"FFFF",X"03E8",X"0000",X"FF01",X"FF00",X"0201",X"03E8",
X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"0224",X"03E8",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"0237",X"03E8",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"0218",X"03E8",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"0060",X"004A",X"000D",X"FFFF",
X"03E8",X"0000",X"FF01",X"FF00",X"0254",X"03E8",X"0006",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"026C",X"03E8",X"0009",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"025C",X"03E8",X"0003",X"00BB",X"0164",X"06DB",X"0276",
X"03E8",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"024E",X"03E8",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"024B",X"03E8",X"0006",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"026A",X"03E8",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0060",X"001D",
X"000E",X"FFFF",X"03E8",X"0000",X"FF01",X"FF00",X"0284",X"03E8",
X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"0286",X"03E8",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"0060",X"0062",X"000F",X"FFFF",X"03E8",
X"0000",X"FF01",X"FF00",X"02DA",X"03E8",X"0009",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"02E5",
X"03E8",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"02E0",
X"03E8",X"0003",X"00BB",X"0164",X"06DB",X"02DF",X"03E8",X"0009",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"02CE",X"03E8",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"02E4",X"03E8",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"02C6",
X"03E8",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"02D7",
X"03E8",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"02C6",X"03E8",X"0007",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0127",X"FF00",X"0060",
X"0035",X"0008",X"FFFF",X"03F2",X"0001",X"FF01",X"FF00",X"0234",
X"03F2",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"020D",X"03F2",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"0234",X"03F2",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"0231",X"03F2",X"0003",X"00BB",X"0164",X"06DB",X"022E",
X"03F2",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"0060",X"0053",X"0009",X"FFFF",
X"03F2",X"0001",X"FF01",X"FF00",X"0256",X"03F2",X"0003",X"00BB",
X"0164",X"06DB",X"0245",X"03F2",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"026B",X"03F2",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0261",X"03F2",X"0003",X"00BB",X"0164",X"06DB",
X"0276",X"03F2",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"025C",X"03F2",X"000A",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
X"0246",X"03F2",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0268",X"03F2",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0060",
X"002C",X"000A",X"FFFF",X"03F2",X"0001",X"FF01",X"FF00",X"0289",
X"03F2",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"029E",X"03F2",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"02BD",X"03F2",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0290",X"03F2",X"0003",
X"00BB",X"0164",X"06DB",X"0060",X"0008",X"000B",X"FFFF",X"03F2",
X"0001",X"FF01",X"FF00",X"0060",X"001C",X"000C",X"FFFF",X"03F2",
X"0001",X"FF01",X"FF00",X"021B",X"03F2",X"0005",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0226",X"03F2",X"0009",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0060",
X"0008",X"000D",X"FFFF",X"03F2",X"0001",X"FF01",X"FF00",X"0060",
X"0022",X"000E",X"FFFF",X"03F2",X"0001",X"FF01",X"FF00",X"0295",
X"03F2",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"0283",X"03F2",X"000A",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"00E0",X"0060",X"0023",X"000F",X"FFFF",X"03F2",X"0001",X"FF01",
X"FF00",X"02C3",X"03F2",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"02D5",X"03F2",X"0003",
X"00BB",X"0164",X"06DB",X"02EE",X"03F2",X"0006",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"01F7",X"FF00",X"0060",X"005F",
X"0008",X"FFFF",X"03FC",X"0002",X"FF01",X"FF00",X"023C",X"03FC",
X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"0204",X"03FC",X"0006",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"0239",X"03FC",X"0005",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0236",X"03FC",X"0007",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0228",X"03FC",X"0006",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0208",X"03FC",
X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"022B",X"03FC",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"020A",X"03FC",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"0226",X"03FC",X"0006",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0060",X"0010",X"0009",
X"FFFF",X"03FC",X"0002",X"FF01",X"FF00",X"027D",X"03FC",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0060",X"0017",X"000A",
X"FFFF",X"03FC",X"0002",X"FF01",X"FF00",X"029F",X"03FC",X"0006",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0297",X"03FC",
X"0003",X"00BB",X"0164",X"06DB",X"0060",X"0049",X"000B",X"FFFF",
X"03FC",X"0002",X"FF01",X"FF00",X"02E3",X"03FC",X"000A",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"00E0",X"02DE",X"03FC",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"02D3",X"03FC",X"0007",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"02F8",X"03FC",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"02CA",X"03FC",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"02F3",X"03FC",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"02E5",
X"03FC",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"006A",X"000C",
X"FFFF",X"03FC",X"0002",X"FF01",X"FF00",X"0234",X"03FC",X"0004",
X"00BB",X"0164",X"06DB",X"0F1B",X"0212",X"03FC",X"0008",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0229",
X"03FC",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"0219",X"03FC",X"000A",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0204",
X"03FC",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"0238",X"03FC",X"0005",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"020F",X"03FC",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"020A",X"03FC",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0209",X"03FC",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0231",
X"03FC",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0060",
X"0046",X"000D",X"FFFF",X"03FC",X"0002",X"FF01",X"FF00",X"0273",
X"03FC",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"024C",X"03FC",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0252",
X"03FC",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"026F",X"03FC",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0275",X"03FC",X"000A",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0276",
X"03FC",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0244",
X"03FC",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"0054",X"000E",
X"FFFF",X"03FC",X"0002",X"FF01",X"FF00",X"028C",X"03FC",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"028A",X"03FC",X"0008",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"02B1",X"03FC",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"02A3",
X"03FC",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"0298",X"03FC",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0280",X"03FC",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0286",X"03FC",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"0291",X"03FC",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"0060",X"0022",X"000F",X"FFFF",X"03FC",X"0002",X"FF01",
X"FF00",X"02DA",X"03FC",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
X"02E8",X"03FC",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"02C4",X"03FC",X"0006",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"0203",X"FF00",X"0060",X"003B",X"0008",
X"FFFF",X"0406",X"0003",X"FF01",X"FF00",X"022C",X"0406",X"0004",
X"00BB",X"0164",X"06DB",X"0F1B",X"0208",X"0406",X"0003",X"00BB",
X"0164",X"06DB",X"0230",X"0406",X"0008",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"021B",X"0406",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0227",X"0406",X"0003",
X"00BB",X"0164",X"06DB",X"023B",X"0406",X"000A",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
X"0060",X"001F",X"0009",X"FFFF",X"0406",X"0003",X"FF01",X"FF00",
X"027C",X"0406",X"0003",X"00BB",X"0164",X"06DB",X"025F",X"0406",
X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"026F",X"0406",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0060",
X"003F",X"000A",X"FFFF",X"0406",X"0003",X"FF01",X"FF00",X"0290",
X"0406",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0297",
X"0406",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"029A",X"0406",X"0009",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"02B3",
X"0406",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"02A2",X"0406",X"0008",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0060",X"0069",
X"000B",X"FFFF",X"0406",X"0003",X"FF01",X"FF00",X"02FF",X"0406",
X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"02F7",X"0406",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"02D1",X"0406",X"0005",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"02CE",X"0406",X"0008",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"02C9",
X"0406",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"02F9",X"0406",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"02D4",X"0406",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"02E8",X"0406",
X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"02C1",X"0406",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"02EC",X"0406",X"0003",X"00BB",X"0164",X"06DB",X"0060",
X"0015",X"000C",X"FFFF",X"0406",X"0003",X"FF01",X"FF00",X"022D",
X"0406",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"0060",X"0010",X"000D",X"FFFF",
X"0406",X"0003",X"FF01",X"FF00",X"0258",X"0406",X"0005",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0060",X"006E",X"000E",X"FFFF",
X"0406",X"0003",X"FF01",X"FF00",X"0297",X"0406",X"0003",X"00BB",
X"0164",X"06DB",X"02A2",X"0406",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"02BC",X"0406",
X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0285",X"0406",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"028A",X"0406",X"000A",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0295",
X"0406",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"029F",X"0406",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"028C",X"0406",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0280",X"0406",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0281",X"0406",
X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"0060",X"006C",X"000F",X"FFFF",X"0406",X"0003",
X"FF01",X"FF00",X"02E2",X"0406",X"0006",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"02F7",X"0406",X"0007",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"02E4",X"0406",X"0009",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"02E0",X"0406",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"02FA",X"0406",X"0004",X"00BB",
X"0164",X"06DB",X"0F1B",X"02E9",X"0406",X"0007",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"02E8",X"0406",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"02C7",
X"0406",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"02DC",X"0406",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"02E3",X"0406",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01A0",X"FF00",
X"0060",X"001A",X"0008",X"FFFF",X"0410",X"0004",X"FF01",X"FF00",
X"0227",X"0410",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"022F",X"0410",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"0060",X"001E",X"0009",X"FFFF",X"0410",X"0004",
X"FF01",X"FF00",X"0265",X"0410",X"0003",X"00BB",X"0164",X"06DB",
X"024F",X"0410",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"024B",X"0410",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0060",X"0008",X"000A",X"FFFF",X"0410",X"0004",X"FF01",X"FF00",
X"0060",X"0025",X"000B",X"FFFF",X"0410",X"0004",X"FF01",X"FF00",
X"02CA",X"0410",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"02F5",
X"0410",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"02F1",X"0410",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0060",X"005E",X"000C",
X"FFFF",X"0410",X"0004",X"FF01",X"FF00",X"021F",X"0410",X"0009",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"021E",X"0410",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
X"023D",X"0410",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"023B",X"0410",X"0005",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"021D",X"0410",X"0005",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0221",X"0410",X"0005",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0214",X"0410",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"0222",X"0410",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0209",
X"0410",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"0060",X"0054",X"000D",X"FFFF",X"0410",
X"0004",X"FF01",X"FF00",X"0279",X"0410",X"0009",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"024B",
X"0410",X"0003",X"00BB",X"0164",X"06DB",X"0240",X"0410",X"0008",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"024A",X"0410",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"024E",X"0410",X"0008",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"026F",X"0410",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0278",X"0410",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0060",
X"006B",X"000E",X"FFFF",X"0410",X"0004",X"FF01",X"FF00",X"02B7",
X"0410",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"02BC",
X"0410",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"02AE",X"0410",X"000A",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"00E0",X"0298",X"0410",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"02B6",X"0410",X"0007",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"0294",X"0410",X"0004",X"00BB",
X"0164",X"06DB",X"0F1B",X"02A1",X"0410",X"0003",X"00BB",X"0164",
X"06DB",X"02B9",X"0410",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0284",X"0410",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"02B4",X"0410",
X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"0060",X"001C",X"000F",X"FFFF",X"0410",X"0004",
X"FF01",X"FF00",X"02DE",X"0410",X"0003",X"00BB",X"0164",X"06DB",
X"02EC",X"0410",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"02F8",
X"0410",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0118",X"FF00",
X"0060",X"0014",X"0008",X"FFFF",X"041A",X"0005",X"FF01",X"FF00",
X"022C",X"041A",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"0060",X"003C",X"0009",X"FFFF",
X"041A",X"0005",X"FF01",X"FF00",X"0247",X"041A",X"0008",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"025F",
X"041A",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"026B",X"041A",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"0255",X"041A",X"0006",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"0256",X"041A",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"0060",X"001E",X"000A",X"FFFF",X"041A",X"0005",X"FF01",X"FF00",
X"0285",X"041A",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"029C",X"041A",X"0006",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0060",X"0019",
X"000B",X"FFFF",X"041A",X"0005",X"FF01",X"FF00",X"02CC",X"041A",
X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"02E7",X"041A",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0060",
X"0054",X"000C",X"FFFF",X"041A",X"0005",X"FF01",X"FF00",X"023F",
X"041A",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"0221",X"041A",X"0006",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0217",X"041A",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"020D",X"041A",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0229",X"041A",
X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"0229",X"041A",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"021E",X"041A",X"0004",X"00BB",
X"0164",X"06DB",X"0F1B",X"0060",X"0017",X"000D",X"FFFF",X"041A",
X"0005",X"FF01",X"FF00",X"0241",X"041A",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"0250",X"041A",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0060",X"001C",X"000E",X"FFFF",X"041A",X"0005",
X"FF01",X"FF00",X"02AA",X"041A",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0296",X"041A",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0060",X"0008",
X"000F",X"FFFF",X"041A",X"0005",X"FF01",X"FF00",X"0181",X"FF00",
X"0060",X"002C",X"0008",X"FFFF",X"0424",X"0006",X"FF01",X"FF00",
X"0222",X"0424",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"021F",X"0424",X"0008",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"021A",
X"0424",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"0060",X"001B",X"0009",X"FFFF",
X"0424",X"0006",X"FF01",X"FF00",X"025D",X"0424",X"0003",X"00BB",
X"0164",X"06DB",X"0269",X"0424",X"000A",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0060",
X"0029",X"000A",X"FFFF",X"0424",X"0006",X"FF01",X"FF00",X"0282",
X"0424",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"02AC",X"0424",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0292",X"0424",
X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"0060",X"005A",X"000B",X"FFFF",X"0424",X"0006",X"FF01",X"FF00",
X"02EB",X"0424",X"0003",X"00BB",X"0164",X"06DB",X"02E1",X"0424",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"02F4",X"0424",X"0005",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"02D7",X"0424",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"02FC",X"0424",X"0003",X"00BB",X"0164",X"06DB",
X"02DD",X"0424",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"02FE",X"0424",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"02E6",X"0424",X"0006",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"02EC",X"0424",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"0060",X"004B",X"000C",X"FFFF",X"0424",X"0006",
X"FF01",X"FF00",X"0234",X"0424",X"0007",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"0218",X"0424",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"0212",X"0424",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0235",X"0424",X"0008",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"020E",X"0424",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"023F",X"0424",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0207",
X"0424",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"0031",X"000D",
X"FFFF",X"0424",X"0006",X"FF01",X"FF00",X"0264",X"0424",X"0003",
X"00BB",X"0164",X"06DB",X"0278",X"0424",X"0007",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0244",X"0424",X"0008",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"0241",X"0424",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"025C",X"0424",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"0025",
X"000E",X"FFFF",X"0424",X"0006",X"FF01",X"FF00",X"02B7",X"0424",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"02B8",X"0424",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"02A2",X"0424",X"0005",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0060",X"0014",X"000F",X"FFFF",X"0424",
X"0006",X"FF01",X"FF00",X"02EB",X"0424",X"0003",X"00BB",X"0164",
X"06DB",X"02DA",X"0424",X"0003",X"00BB",X"0164",X"06DB",X"027F",
X"FF00",X"0060",X"0063",X"0008",X"FFFF",X"042E",X"0007",X"FF01",
X"FF00",X"0238",X"042E",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"0222",X"042E",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"021C",X"042E",
X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"023E",X"042E",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"0219",X"042E",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"022E",X"042E",
X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0204",X"042E",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"023C",X"042E",X"0006",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"023B",X"042E",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0205",X"042E",
X"0003",X"00BB",X"0164",X"06DB",X"0060",X"005D",X"0009",X"FFFF",
X"042E",X"0007",X"FF01",X"FF00",X"026A",X"042E",X"0008",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"027D",
X"042E",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"027E",X"042E",
X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"0278",X"042E",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0251",X"042E",X"0003",X"00BB",X"0164",X"06DB",
X"0244",X"042E",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"0251",X"042E",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"0246",X"042E",X"000A",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"00E0",X"0253",X"042E",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0060",X"005C",X"000A",X"FFFF",X"042E",X"0007",X"FF01",
X"FF00",X"0282",X"042E",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0287",X"042E",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"0298",X"042E",X"000A",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
X"0287",X"042E",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"02B5",X"042E",X"0003",X"00BB",
X"0164",X"06DB",X"029D",X"042E",X"0007",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"02B8",X"042E",X"0008",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0283",
X"042E",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"0039",X"000B",
X"FFFF",X"042E",X"0007",X"FF01",X"FF00",X"02CD",X"042E",X"0003",
X"00BB",X"0164",X"06DB",X"02C2",X"042E",X"000A",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
X"02D6",X"042E",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"02E6",
X"042E",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"02FE",X"042E",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"02CF",X"042E",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"002F",
X"000C",X"FFFF",X"042E",X"0007",X"FF01",X"FF00",X"021F",X"042E",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"022B",
X"042E",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0234",
X"042E",X"0003",X"00BB",X"0164",X"06DB",X"0211",X"042E",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0214",
X"042E",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"005B",X"000D",
X"FFFF",X"042E",X"0007",X"FF01",X"FF00",X"024C",X"042E",X"0004",
X"00BB",X"0164",X"06DB",X"0F1B",X"025A",X"042E",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"0266",X"042E",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"0257",X"042E",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0265",X"042E",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"027B",X"042E",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0245",X"042E",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"026C",X"042E",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0250",X"042E",
X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"0060",X"0069",X"000E",X"FFFF",X"042E",X"0007",X"FF01",X"FF00",
X"0295",X"042E",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"02BA",X"042E",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"02AA",X"042E",X"0005",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0291",X"042E",X"0006",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0283",X"042E",X"0006",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"02A0",X"042E",
X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"02AE",X"042E",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0297",X"042E",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"029D",X"042E",
X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"02B7",X"042E",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"0060",X"0035",X"000F",X"FFFF",X"042E",X"0007",X"FF01",
X"FF00",X"02C9",X"042E",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"02F3",X"042E",X"000A",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"00E0",X"02FB",X"042E",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"02FD",X"042E",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"01CB",X"FF00",
X"0060",X"0040",X"0008",X"FFFF",X"0438",X"0008",X"FF01",X"FF00",
X"0233",X"0438",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"0220",X"0438",X"0009",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0214",
X"0438",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"020D",X"0438",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0212",X"0438",
X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"0060",X"005C",X"0009",X"FFFF",X"0438",X"0008",X"FF01",X"FF00",
X"0241",X"0438",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0263",X"0438",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0260",
X"0438",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"0261",X"0438",X"0007",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0264",X"0438",X"0003",
X"00BB",X"0164",X"06DB",X"024E",X"0438",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"0265",X"0438",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"025E",X"0438",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
X"024E",X"0438",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"0060",X"0021",X"000A",X"FFFF",
X"0438",X"0008",X"FF01",X"FF00",X"02A5",X"0438",X"0008",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"02B3",
X"0438",X"0003",X"00BB",X"0164",X"06DB",X"028E",X"0438",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0060",X"0021",X"000B",
X"FFFF",X"0438",X"0008",X"FF01",X"FF00",X"02C7",X"0438",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"02DC",X"0438",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"02CB",
X"0438",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0060",X"0061",
X"000C",X"FFFF",X"0438",X"0008",X"FF01",X"FF00",X"0231",X"0438",
X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"023F",X"0438",X"0008",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0236",X"0438",X"0003",
X"00BB",X"0164",X"06DB",X"021E",X"0438",X"000A",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
X"0210",X"0438",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"022A",X"0438",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"0219",X"0438",X"0008",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0235",X"0438",
X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"0218",X"0438",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0060",
X"005F",X"000D",X"FFFF",X"0438",X"0008",X"FF01",X"FF00",X"026E",
X"0438",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"025C",X"0438",X"0005",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"025D",X"0438",X"0008",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0242",
X"0438",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"024D",X"0438",
X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"025F",X"0438",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0245",X"0438",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"0262",X"0438",X"0009",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"025F",
X"0438",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0060",X"0008",
X"000E",X"FFFF",X"0438",X"0008",X"FF01",X"FF00",X"0060",X"0023",
X"000F",X"FFFF",X"0438",X"0008",X"FF01",X"FF00",X"02F4",X"0438",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"02EB",
X"0438",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"02C9",X"0438",X"0003",X"00BB",X"0164",
X"06DB",X"018C",X"FF00",X"0060",X"0012",X"0008",X"FFFF",X"0442",
X"0009",X"FF01",X"FF00",X"0205",X"0442",X"0007",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0060",X"0046",X"0009",
X"FFFF",X"0442",X"0009",X"FF01",X"FF00",X"024D",X"0442",X"0008",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"024D",X"0442",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0258",X"0442",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"0259",X"0442",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0257",X"0442",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"0060",X"0043",X"000A",X"FFFF",X"0442",
X"0009",X"FF01",X"FF00",X"0295",X"0442",X"0009",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0291",
X"0442",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0296",
X"0442",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"0289",X"0442",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"02A3",
X"0442",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"02BF",X"0442",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0060",X"002A",
X"000B",X"FFFF",X"0442",X"0009",X"FF01",X"FF00",X"02E7",X"0442",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"02C6",
X"0442",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"02E5",X"0442",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"02E1",X"0442",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0060",X"0026",X"000C",X"FFFF",X"0442",X"0009",X"FF01",X"FF00",
X"0209",X"0442",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0227",
X"0442",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"0238",X"0442",X"0003",X"00BB",X"0164",X"06DB",X"020B",X"0442",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0060",X"0054",
X"000D",X"FFFF",X"0442",X"0009",X"FF01",X"FF00",X"0250",X"0442",
X"0003",X"00BB",X"0164",X"06DB",X"0279",X"0442",X"000A",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"00E0",X"025F",X"0442",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"024E",X"0442",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"025D",X"0442",X"0008",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"027C",X"0442",X"0008",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"0251",X"0442",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"025E",X"0442",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"0060",X"0043",X"000E",X"FFFF",X"0442",X"0009",
X"FF01",X"FF00",X"0293",X"0442",X"000A",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0291",
X"0442",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"0284",X"0442",X"0005",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0297",X"0442",X"0005",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"02AF",X"0442",X"0008",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0291",X"0442",
X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0060",X"0008",X"000F",
X"FFFF",X"0442",X"0009",X"FF01",X"FF00",X"01DF",X"FF00",X"0060",
X"0038",X"0008",X"FFFF",X"044C",X"000A",X"FF01",X"FF00",X"0222",
X"044C",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"022F",X"044C",X"0003",X"00BB",X"0164",X"06DB",X"0238",
X"044C",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"022C",X"044C",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"020C",
X"044C",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0220",X"044C",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0060",
X"002A",X"0009",X"FFFF",X"044C",X"000A",X"FF01",X"FF00",X"026B",
X"044C",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"024D",X"044C",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"0258",X"044C",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"024C",X"044C",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0060",X"0029",X"000A",X"FFFF",X"044C",X"000A",X"FF01",
X"FF00",X"029E",X"044C",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"02AE",X"044C",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"029F",X"044C",X"0003",X"00BB",
X"0164",X"06DB",X"0293",X"044C",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0060",X"0054",X"000B",X"FFFF",X"044C",X"000A",
X"FF01",X"FF00",X"02EB",X"044C",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"02D7",X"044C",
X"0003",X"00BB",X"0164",X"06DB",X"02C8",X"044C",X"0004",X"00BB",
X"0164",X"06DB",X"0F1B",X"02D5",X"044C",X"0008",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"02F8",X"044C",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"02DC",
X"044C",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"02E3",X"044C",X"0003",X"00BB",X"0164",
X"06DB",X"02D4",X"044C",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0060",X"0008",
X"000C",X"FFFF",X"044C",X"000A",X"FF01",X"FF00",X"0060",X"003A",
X"000D",X"FFFF",X"044C",X"000A",X"FF01",X"FF00",X"0271",X"044C",
X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"0277",X"044C",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"0277",X"044C",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0246",X"044C",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"024D",X"044C",X"0003",X"00BB",X"0164",X"06DB",
X"0060",X"005B",X"000E",X"FFFF",X"044C",X"000A",X"FF01",X"FF00",
X"029D",X"044C",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"02B9",X"044C",X"0003",X"00BB",X"0164",X"06DB",X"02AD",
X"044C",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"02AA",X"044C",
X"0003",X"00BB",X"0164",X"06DB",X"0281",X"044C",X"000A",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"00E0",X"0291",X"044C",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0286",X"044C",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0291",
X"044C",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"02A4",X"044C",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"0060",X"0061",X"000F",X"FFFF",X"044C",
X"000A",X"FF01",X"FF00",X"02CE",X"044C",X"0009",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"02F3",
X"044C",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"02E8",X"044C",X"0009",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"02D3",
X"044C",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"02C3",X"044C",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"02C5",X"044C",X"0006",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"02D8",X"044C",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"02D6",X"044C",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"01DA",X"FF00",X"0060",X"0026",
X"0008",X"FFFF",X"0456",X"000B",X"FF01",X"FF00",X"0227",X"0456",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0209",
X"0456",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"020B",X"0456",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"0060",X"004E",X"0009",X"FFFF",
X"0456",X"000B",X"FF01",X"FF00",X"0268",X"0456",X"0008",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0260",
X"0456",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0270",X"0456",
X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"026F",X"0456",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"024C",X"0456",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0242",X"0456",
X"0003",X"00BB",X"0164",X"06DB",X"024B",X"0456",X"0005",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0264",X"0456",X"0003",X"00BB",
X"0164",X"06DB",X"0060",X"0052",X"000A",X"FFFF",X"0456",X"000B",
X"FF01",X"FF00",X"0287",X"0456",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0282",X"0456",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"02B2",X"0456",X"0008",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"02AB",X"0456",X"0006",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"02B8",X"0456",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"0285",X"0456",X"0003",X"00BB",X"0164",
X"06DB",X"0297",X"0456",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"02B3",X"0456",X"0006",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"0060",X"0011",X"000B",X"FFFF",
X"0456",X"000B",X"FF01",X"FF00",X"02F0",X"0456",X"0006",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0060",X"002A",X"000C",
X"FFFF",X"0456",X"000B",X"FF01",X"FF00",X"020F",X"0456",X"0009",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"0234",X"0456",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"0221",X"0456",X"0008",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0060",
X"002D",X"000D",X"FFFF",X"0456",X"000B",X"FF01",X"FF00",X"0242",
X"0456",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"0246",X"0456",X"0003",X"00BB",
X"0164",X"06DB",X"026D",X"0456",X"0008",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0267",X"0456",X"0004",
X"00BB",X"0164",X"06DB",X"0F1B",X"0060",X"0058",X"000E",X"FFFF",
X"0456",X"000B",X"FF01",X"FF00",X"02B8",X"0456",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"0285",X"0456",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0290",
X"0456",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"02A8",X"0456",X"000A",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
X"02A0",X"0456",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"02A9",X"0456",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"02AD",X"0456",X"0006",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"02B4",X"0456",X"0004",
X"00BB",X"0164",X"06DB",X"0F1B",X"0060",X"0052",X"000F",X"FFFF",
X"0456",X"000B",X"FF01",X"FF00",X"02C4",X"0456",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"02EE",X"0456",
X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"02E3",X"0456",X"0003",
X"00BB",X"0164",X"06DB",X"02FD",X"0456",X"0009",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"02D0",
X"0456",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"02EF",X"0456",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"02C2",X"0456",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"02DA",X"0456",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980");

Constant LinkDat2_Size : Integer := 5291;
Type LinkDat2_Array is Array(0 to LinkDat2_Size - 1) of std_logic_vector(15 downto 0);
Constant LinkDat2 : LinkDat2_Array := 
(X"01E8",X"01D7",X"FF00",X"0060",X"004C",X"0010",X"FFFF",X"03E8",X"0000",
X"FF01",X"FF00",X"042F",X"03E8",X"0007",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"0430",X"03E8",X"0004",X"00BB",
X"0164",X"06DB",X"0F1B",X"040E",X"03E8",X"0003",X"00BB",X"0164",
X"06DB",X"0423",X"03E8",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"0438",X"03E8",X"000A",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"00E0",X"0425",X"03E8",X"0003",X"00BB",X"0164",X"06DB",X"041C",
X"03E8",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"043A",X"03E8",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"000E",
X"0011",X"FFFF",X"03E8",X"0000",X"FF01",X"FF00",X"0444",X"03E8",
X"0003",X"00BB",X"0164",X"06DB",X"0060",X"004E",X"0012",X"FFFF",
X"03E8",X"0000",X"FF01",X"FF00",X"048E",X"03E8",X"0004",X"00BB",
X"0164",X"06DB",X"0F1B",X"04B5",X"03E8",X"0008",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"04BA",X"03E8",
X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"0488",X"03E8",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0495",X"03E8",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"04A1",X"03E8",
X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"04B6",X"03E8",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"0060",X"0034",X"0013",X"FFFF",X"03E8",X"0000",
X"FF01",X"FF00",X"04E0",X"03E8",X"0008",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"04E5",X"03E8",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"04E4",
X"03E8",X"0003",X"00BB",X"0164",X"06DB",X"04E4",X"03E8",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"04D3",
X"03E8",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0060",X"0014",
X"0014",X"FFFF",X"03E8",X"0000",X"FF01",X"FF00",X"0421",X"03E8",
X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"0060",X"004A",X"0015",X"FFFF",X"03E8",X"0000",
X"FF01",X"FF00",X"0444",X"03E8",X"0007",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"0454",X"03E8",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"044E",X"03E8",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"045C",X"03E8",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0458",X"03E8",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0473",
X"03E8",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"0060",X"0030",X"0016",X"FFFF",
X"03E8",X"0000",X"FF01",X"FF00",X"049E",X"03E8",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"0486",X"03E8",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"048A",
X"03E8",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"049F",X"03E8",X"0007",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"0060",X"006B",X"0017",X"FFFF",
X"03E8",X"0000",X"FF01",X"FF00",X"04FF",X"03E8",X"0006",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"04D7",X"03E8",X"0008",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"04F0",X"03E8",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"04EE",X"03E8",X"0006",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"04C9",X"03E8",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"04ED",X"03E8",X"0006",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"04CE",X"03E8",X"0003",X"00BB",X"0164",
X"06DB",X"04E0",X"03E8",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"04D3",X"03E8",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"04DA",X"03E8",X"0009",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0249",
X"FF00",X"0060",X"0059",X"0010",X"FFFF",X"03F2",X"0001",X"FF01",
X"FF00",X"042C",X"03F2",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"0436",X"03F2",X"0009",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"0437",X"03F2",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"0420",X"03F2",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"040A",X"03F2",
X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"0433",X"03F2",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"0417",X"03F2",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0437",X"03F2",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"0060",X"0067",X"0011",X"FFFF",X"03F2",X"0001",
X"FF01",X"FF00",X"045F",X"03F2",X"0006",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"045A",X"03F2",X"0008",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0472",X"03F2",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"044C",
X"03F2",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"0462",X"03F2",X"0003",X"00BB",
X"0164",X"06DB",X"0454",X"03F2",X"0007",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"0479",X"03F2",X"000A",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"00E0",X"044C",X"03F2",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"047B",X"03F2",
X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"0060",X"0011",X"0012",X"FFFF",X"03F2",X"0001",X"FF01",
X"FF00",X"0494",X"03F2",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"0060",X"0065",X"0013",X"FFFF",X"03F2",X"0001",
X"FF01",X"FF00",X"04C2",X"03F2",X"0008",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"04FC",X"03F2",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"04EC",X"03F2",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"04D0",X"03F2",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"04C7",X"03F2",X"000A",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"04E0",
X"03F2",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"04C7",X"03F2",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"04D7",X"03F2",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"04D6",
X"03F2",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0060",
X"0075",X"0014",X"FFFF",X"03F2",X"0001",X"FF01",X"FF00",X"041D",
X"03F2",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"0418",X"03F2",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"0408",X"03F2",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0428",X"03F2",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0425",
X"03F2",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"0428",X"03F2",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0430",X"03F2",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
X"0405",X"03F2",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"043D",X"03F2",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"0406",X"03F2",X"0007",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"0060",X"0036",X"0015",X"FFFF",
X"03F2",X"0001",X"FF01",X"FF00",X"0466",X"03F2",X"0004",X"00BB",
X"0164",X"06DB",X"0F1B",X"0469",X"03F2",X"0005",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"047C",X"03F2",X"0003",X"00BB",X"0164",
X"06DB",X"0471",X"03F2",X"0003",X"00BB",X"0164",X"06DB",X"0445",
X"03F2",X"0003",X"00BB",X"0164",X"06DB",X"0473",X"03F2",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"0060",X"003A",X"0016",X"FFFF",X"03F2",X"0001",
X"FF01",X"FF00",X"04AE",X"03F2",X"000A",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0495",
X"03F2",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"04B4",X"03F2",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"04BA",X"03F2",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"0488",X"03F2",X"0007",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"0060",X"002C",X"0017",X"FFFF",
X"03F2",X"0001",X"FF01",X"FF00",X"04E1",X"03F2",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"04E5",X"03F2",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"04D8",X"03F2",X"000A",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
X"01F4",X"FF00",X"0060",X"0051",X"0010",X"FFFF",X"03FC",X"0002",
X"FF01",X"FF00",X"0411",X"03FC",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0413",X"03FC",
X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"0411",X"03FC",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"0413",X"03FC",X"0003",X"00BB",X"0164",X"06DB",
X"042A",X"03FC",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"0417",X"03FC",X"0004",X"00BB",
X"0164",X"06DB",X"0F1B",X"0400",X"03FC",X"0007",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0422",X"03FC",X"0003",
X"00BB",X"0164",X"06DB",X"0060",X"004A",X"0011",X"FFFF",X"03FC",
X"0002",X"FF01",X"FF00",X"0469",X"03FC",X"0008",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"046E",X"03FC",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"0470",X"03FC",X"000A",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
X"0467",X"03FC",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"0470",X"03FC",X"0003",X"00BB",X"0164",X"06DB",
X"0457",X"03FC",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0060",X"002A",X"0012",
X"FFFF",X"03FC",X"0002",X"FF01",X"FF00",X"04B1",X"03FC",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0493",
X"03FC",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"04A0",X"03FC",X"000A",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0060",
X"0046",X"0013",X"FFFF",X"03FC",X"0002",X"FF01",X"FF00",X"04E9",
X"03FC",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"04EB",
X"03FC",X"0003",X"00BB",X"0164",X"06DB",X"04C1",X"03FC",X"0003",
X"00BB",X"0164",X"06DB",X"04DF",X"03FC",X"0006",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"04C6",X"03FC",X"0004",X"00BB",
X"0164",X"06DB",X"0F1B",X"04DF",X"03FC",X"0005",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"04F8",X"03FC",X"0009",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"04F9",
X"03FC",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"0022",X"0014",
X"FFFF",X"03FC",X"0002",X"FF01",X"FF00",X"0416",X"03FC",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0417",X"03FC",X"0006",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"040D",X"03FC",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0060",
X"004A",X"0015",X"FFFF",X"03FC",X"0002",X"FF01",X"FF00",X"046F",
X"03FC",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"047F",X"03FC",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"045B",X"03FC",X"0003",X"00BB",X"0164",X"06DB",
X"044F",X"03FC",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"0449",X"03FC",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"0467",X"03FC",X"0006",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"0447",X"03FC",X"0003",X"00BB",X"0164",
X"06DB",X"0444",X"03FC",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0060",X"001F",X"0016",X"FFFF",X"03FC",X"0002",X"FF01",
X"FF00",X"04A2",X"03FC",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"0484",X"03FC",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"0482",X"03FC",X"0003",X"00BB",X"0164",X"06DB",
X"0060",X"005C",X"0017",X"FFFF",X"03FC",X"0002",X"FF01",X"FF00",
X"04D2",X"03FC",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"04DA",X"03FC",X"0008",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"04D9",
X"03FC",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"04C4",
X"03FC",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"04C8",X"03FC",X"0003",X"00BB",X"0164",
X"06DB",X"04DF",X"03FC",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"04D2",X"03FC",X"0007",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"04D3",X"03FC",X"0003",
X"00BB",X"0164",X"06DB",X"04D7",X"03FC",X"0006",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"01C1",X"FF00",X"0060",X"0064",
X"0010",X"FFFF",X"0406",X"0003",X"FF01",X"FF00",X"043F",X"0406",
X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"0412",X"0406",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"043E",X"0406",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"0430",X"0406",X"0007",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0432",X"0406",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0407",
X"0406",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"0412",X"0406",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"043C",X"0406",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"043B",X"0406",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0060",X"0028",X"0011",X"FFFF",X"0406",X"0003",
X"FF01",X"FF00",X"0446",X"0406",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"044C",X"0406",X"000A",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0471",
X"0406",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"0060",X"005C",X"0012",X"FFFF",X"0406",X"0003",
X"FF01",X"FF00",X"04A7",X"0406",X"0007",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"04B1",X"0406",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"04AE",X"0406",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0482",X"0406",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"0494",X"0406",X"000A",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"04A5",
X"0406",X"0003",X"00BB",X"0164",X"06DB",X"0494",X"0406",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"0494",X"0406",X"0003",X"00BB",X"0164",X"06DB",
X"049E",X"0406",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"0029",
X"0013",X"FFFF",X"0406",X"0003",X"FF01",X"FF00",X"04FE",X"0406",
X"0003",X"00BB",X"0164",X"06DB",X"04D9",X"0406",X"0003",X"00BB",
X"0164",X"06DB",X"04DF",X"0406",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"04F4",X"0406",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0060",
X"0008",X"0014",X"FFFF",X"0406",X"0003",X"FF01",X"FF00",X"0060",
X"0024",X"0015",X"FFFF",X"0406",X"0003",X"FF01",X"FF00",X"0448",
X"0406",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"046F",
X"0406",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"0450",X"0406",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"0060",X"0033",X"0016",X"FFFF",X"0406",
X"0003",X"FF01",X"FF00",X"048C",X"0406",X"0006",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"049B",X"0406",X"0008",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"04A6",
X"0406",X"0003",X"00BB",X"0164",X"06DB",X"04BF",X"0406",X"0004",
X"00BB",X"0164",X"06DB",X"0F1B",X"048F",X"0406",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0060",X"004F",
X"0017",X"FFFF",X"0406",X"0003",X"FF01",X"FF00",X"04C6",X"0406",
X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"04EB",X"0406",X"0003",X"00BB",X"0164",X"06DB",X"04E4",X"0406",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"04FB",
X"0406",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"04D8",X"0406",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"04F0",X"0406",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
X"04DF",X"0406",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"04FA",X"0406",X"0006",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0181",X"FF00",X"0060",
X"0043",X"0010",X"FFFF",X"0410",X"0004",X"FF01",X"FF00",X"0423",
X"0410",X"0003",X"00BB",X"0164",X"06DB",X"0405",X"0410",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"043F",X"0410",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"040B",X"0410",X"0006",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"0424",X"0410",X"0007",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0417",X"0410",X"0003",
X"00BB",X"0164",X"06DB",X"042F",X"0410",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"0060",X"003E",X"0011",X"FFFF",X"0410",X"0004",
X"FF01",X"FF00",X"0478",X"0410",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"0441",X"0410",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
X"044E",X"0410",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"046F",X"0410",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"0466",X"0410",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"046F",X"0410",X"0003",X"00BB",X"0164",X"06DB",
X"0060",X"0008",X"0012",X"FFFF",X"0410",X"0004",X"FF01",X"FF00",
X"0060",X"005E",X"0013",X"FFFF",X"0410",X"0004",X"FF01",X"FF00",
X"04E5",X"0410",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"04D9",X"0410",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"04C4",X"0410",X"0003",X"00BB",X"0164",X"06DB",X"04FF",X"0410",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"04FC",
X"0410",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"04DD",X"0410",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
X"04D6",X"0410",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"04CC",X"0410",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"04E2",X"0410",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0060",X"000F",
X"0014",X"FFFF",X"0410",X"0004",X"FF01",X"FF00",X"040F",X"0410",
X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0060",X"0025",X"0015",
X"FFFF",X"0410",X"0004",X"FF01",X"FF00",X"0442",X"0410",X"0003",
X"00BB",X"0164",X"06DB",X"044A",X"0410",X"0006",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"0456",X"0410",X"0005",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0446",X"0410",X"0003",X"00BB",
X"0164",X"06DB",X"0060",X"0012",X"0016",X"FFFF",X"0410",X"0004",
X"FF01",X"FF00",X"049F",X"0410",X"0007",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"0060",X"0052",X"0017",X"FFFF",
X"0410",X"0004",X"FF01",X"FF00",X"04F5",X"0410",X"000A",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"00E0",X"04C5",X"0410",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"04C0",X"0410",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"04E8",X"0410",X"0008",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"04DE",X"0410",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"04F5",X"0410",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"04F6",X"0410",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"01BB",X"FF00",
X"0060",X"004B",X"0010",X"FFFF",X"041A",X"0005",X"FF01",X"FF00",
X"0431",X"041A",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"042B",X"041A",X"0008",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"041F",X"041A",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0404",X"041A",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0431",X"041A",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0418",
X"041A",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"042C",X"041A",X"0005",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0060",X"001B",X"0011",X"FFFF",X"041A",
X"0005",X"FF01",X"FF00",X"045C",X"041A",X"0006",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"0479",X"041A",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0060",X"001A",
X"0012",X"FFFF",X"041A",X"0005",X"FF01",X"FF00",X"0485",X"041A",
X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0484",X"041A",X"0008",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"0060",X"0066",X"0013",X"FFFF",X"041A",X"0005",X"FF01",X"FF00",
X"04FD",X"041A",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"04DF",X"041A",X"000A",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
X"04DB",X"041A",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"04FF",X"041A",X"0006",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"04E7",X"041A",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"04D6",X"041A",X"0007",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"04E1",X"041A",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"04D3",X"041A",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0060",X"0033",
X"0014",X"FFFF",X"041A",X"0005",X"FF01",X"FF00",X"0405",X"041A",
X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0428",X"041A",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0408",
X"041A",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"0436",X"041A",X"0003",X"00BB",X"0164",X"06DB",
X"0412",X"041A",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"0060",X"0060",X"0015",X"FFFF",X"041A",X"0005",X"FF01",
X"FF00",X"0453",X"041A",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0456",X"041A",
X"0003",X"00BB",X"0164",X"06DB",X"0445",X"041A",X"0005",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0442",X"041A",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"046D",X"041A",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"0466",X"041A",X"0006",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0471",X"041A",X"0009",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"0473",X"041A",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"0467",X"041A",X"0003",X"00BB",X"0164",
X"06DB",X"0060",X"0038",X"0016",X"FFFF",X"041A",X"0005",X"FF01",
X"FF00",X"0498",X"041A",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
X"04AF",X"041A",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"0491",X"041A",X"0008",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0494",
X"041A",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"0489",X"041A",X"0003",X"00BB",X"0164",
X"06DB",X"0060",X"0008",X"0017",X"FFFF",X"041A",X"0005",X"FF01",
X"FF00",X"01EA",X"FF00",X"0060",X"0053",X"0010",X"FFFF",X"0424",
X"0006",X"FF01",X"FF00",X"041E",X"0424",X"0007",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0438",X"0424",X"0008",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"041A",X"0424",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"0417",X"0424",X"0009",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0432",
X"0424",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"0400",X"0424",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"040F",X"0424",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0060",X"003E",
X"0011",X"FFFF",X"0424",X"0006",X"FF01",X"FF00",X"0458",X"0424",
X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0450",X"0424",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0462",
X"0424",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0478",X"0424",
X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"045A",X"0424",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
X"0477",X"0424",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"0060",X"004B",X"0012",X"FFFF",
X"0424",X"0006",X"FF01",X"FF00",X"049F",X"0424",X"000A",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"00E0",X"04A7",X"0424",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"0495",X"0424",X"0004",
X"00BB",X"0164",X"06DB",X"0F1B",X"0489",X"0424",X"0004",X"00BB",
X"0164",X"06DB",X"0F1B",X"04A8",X"0424",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"04A3",X"0424",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"048D",X"0424",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"04B1",X"0424",X"0003",X"00BB",X"0164",X"06DB",X"0060",
X"0039",X"0013",X"FFFF",X"0424",X"0006",X"FF01",X"FF00",X"04FE",
X"0424",X"0003",X"00BB",X"0164",X"06DB",X"04F6",X"0424",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"04D4",X"0424",X"0003",
X"00BB",X"0164",X"06DB",X"04C3",X"0424",X"0009",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"04FD",
X"0424",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"04D7",X"0424",
X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"0060",X"004F",X"0014",X"FFFF",X"0424",X"0006",X"FF01",X"FF00",
X"042D",X"0424",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"043F",X"0424",X"0003",X"00BB",X"0164",
X"06DB",X"042B",X"0424",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"043E",X"0424",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"0414",X"0424",X"0006",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"0428",X"0424",X"0008",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"041A",
X"0424",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0419",X"0424",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0060",
X"0018",X"0015",X"FFFF",X"0424",X"0006",X"FF01",X"FF00",X"045F",
X"0424",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"0443",X"0424",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0060",
X"001E",X"0016",X"FFFF",X"0424",X"0006",X"FF01",X"FF00",X"04A9",
X"0424",X"0003",X"00BB",X"0164",X"06DB",X"048E",X"0424",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"04A9",
X"0424",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"004E",X"0017",
X"FFFF",X"0424",X"0006",X"FF01",X"FF00",X"04EE",X"0424",X"0003",
X"00BB",X"0164",X"06DB",X"04CB",X"0424",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"04F4",X"0424",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"04E9",X"0424",
X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"04FD",X"0424",X"0004",
X"00BB",X"0164",X"06DB",X"0F1B",X"04ED",X"0424",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"04E0",X"0424",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"04F7",X"0424",X"0005",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"01D8",X"FF00",X"0060",X"0061",X"0010",
X"FFFF",X"042E",X"0007",X"FF01",X"FF00",X"042D",X"042E",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"040A",
X"042E",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0434",X"042E",
X"0003",X"00BB",X"0164",X"06DB",X"0424",X"042E",X"0006",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0420",X"042E",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"043B",X"042E",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0438",X"042E",X"0008",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"043F",X"042E",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"042D",X"042E",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"0060",X"001E",
X"0011",X"FFFF",X"042E",X"0007",X"FF01",X"FF00",X"047D",X"042E",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"047C",X"042E",X"0006",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"0060",X"004F",X"0012",X"FFFF",
X"042E",X"0007",X"FF01",X"FF00",X"0494",X"042E",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"0484",X"042E",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"049E",X"042E",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"0496",X"042E",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"04B8",X"042E",
X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"04B4",X"042E",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"04A5",X"042E",X"0006",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"0060",X"000E",X"0013",X"FFFF",X"042E",
X"0007",X"FF01",X"FF00",X"04F8",X"042E",X"0003",X"00BB",X"0164",
X"06DB",X"0060",X"0047",X"0014",X"FFFF",X"042E",X"0007",X"FF01",
X"FF00",X"0417",X"042E",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0418",X"042E",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"0414",X"042E",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"0400",X"042E",X"0003",X"00BB",X"0164",X"06DB",
X"0423",X"042E",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0403",X"042E",X"0006",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"042C",X"042E",
X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"0060",X"0066",X"0015",X"FFFF",X"042E",X"0007",X"FF01",X"FF00",
X"0461",X"042E",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0457",
X"042E",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"0442",X"042E",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0455",X"042E",
X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0466",X"042E",X"0004",
X"00BB",X"0164",X"06DB",X"0F1B",X"0479",X"042E",X"0003",X"00BB",
X"0164",X"06DB",X"044F",X"042E",X"0009",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"047D",X"042E",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"0476",X"042E",X"0007",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"047B",X"042E",X"0006",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0060",X"0028",
X"0016",X"FFFF",X"042E",X"0007",X"FF01",X"FF00",X"0480",X"042E",
X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"0489",X"042E",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"04AF",X"042E",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0060",X"0025",
X"0017",X"FFFF",X"042E",X"0007",X"FF01",X"FF00",X"04F7",X"042E",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"04E4",
X"042E",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"04CB",X"042E",X"0004",X"00BB",
X"0164",X"06DB",X"0F1B",X"0112",X"FF00",X"0060",X"0013",X"0010",
X"FFFF",X"0438",X"0008",X"FF01",X"FF00",X"040B",X"0438",X"0008",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"0060",X"0008",X"0011",X"FFFF",X"0438",X"0008",X"FF01",X"FF00",
X"0060",X"0032",X"0012",X"FFFF",X"0438",X"0008",X"FF01",X"FF00",
X"04AA",X"0438",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"048A",X"0438",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"04AA",X"0438",X"0003",X"00BB",X"0164",X"06DB",X"0495",
X"0438",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"04B5",X"0438",X"0003",X"00BB",
X"0164",X"06DB",X"0060",X"001E",X"0013",X"FFFF",X"0438",X"0008",
X"FF01",X"FF00",X"04DD",X"0438",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"04FA",X"0438",X"0003",X"00BB",X"0164",X"06DB",X"04F8",
X"0438",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"0060",X"0027",X"0014",X"FFFF",X"0438",X"0008",X"FF01",X"FF00",
X"0412",X"0438",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0407",X"0438",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"043D",X"0438",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0060",
X"0031",X"0015",X"FFFF",X"0438",X"0008",X"FF01",X"FF00",X"047E",
X"0438",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"0462",X"0438",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"045B",X"0438",X"0004",
X"00BB",X"0164",X"06DB",X"0F1B",X"047F",X"0438",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"0060",X"0022",X"0016",X"FFFF",X"0438",X"0008",X"FF01",X"FF00",
X"048B",X"0438",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"04AA",X"0438",X"0003",
X"00BB",X"0164",X"06DB",X"0491",X"0438",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"0060",X"002B",X"0017",X"FFFF",X"0438",X"0008",
X"FF01",X"FF00",X"04CB",X"0438",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"04D9",X"0438",X"0003",X"00BB",X"0164",X"06DB",
X"04C2",X"0438",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"04E6",X"0438",X"0006",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"018D",X"FF00",X"0060",
X"000E",X"0010",X"FFFF",X"0442",X"0009",X"FF01",X"FF00",X"0404",
X"0442",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"0039",X"0011",
X"FFFF",X"0442",X"0009",X"FF01",X"FF00",X"045F",X"0442",X"000A",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"00E0",X"044C",X"0442",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"0473",X"0442",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0461",X"0442",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"0463",X"0442",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0060",X"004A",
X"0012",X"FFFF",X"0442",X"0009",X"FF01",X"FF00",X"04B6",X"0442",
X"0003",X"00BB",X"0164",X"06DB",X"049B",X"0442",X"0003",X"00BB",
X"0164",X"06DB",X"0483",X"0442",X"0003",X"00BB",X"0164",X"06DB",
X"0490",X"0442",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"04A2",X"0442",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"049F",X"0442",X"0004",X"00BB",
X"0164",X"06DB",X"0F1B",X"048A",X"0442",X"000A",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
X"0496",X"0442",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0060",X"0032",X"0013",X"FFFF",X"0442",X"0009",X"FF01",X"FF00",
X"04C7",X"0442",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"04E4",X"0442",X"0003",X"00BB",X"0164",X"06DB",X"04EA",X"0442",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"04F4",
X"0442",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"04D2",X"0442",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"0060",X"0030",X"0014",X"FFFF",X"0442",X"0009",
X"FF01",X"FF00",X"0428",X"0442",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"0433",X"0442",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"041E",X"0442",X"0003",X"00BB",X"0164",X"06DB",
X"041F",X"0442",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"0416",X"0442",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"0060",X"0008",X"0015",X"FFFF",X"0442",X"0009",
X"FF01",X"FF00",X"0060",X"004C",X"0016",X"FFFF",X"0442",X"0009",
X"FF01",X"FF00",X"0496",X"0442",X"000A",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0484",
X"0442",X"0003",X"00BB",X"0164",X"06DB",X"04A4",X"0442",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"04A5",X"0442",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0488",X"0442",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"04B4",X"0442",X"0004",
X"00BB",X"0164",X"06DB",X"0F1B",X"04A7",X"0442",X"0009",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"04A6",X"0442",X"0003",X"00BB",X"0164",X"06DB",X"0060",X"0044",
X"0017",X"FFFF",X"0442",X"0009",X"FF01",X"FF00",X"04EB",X"0442",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"04F2",X"0442",
X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"04DA",X"0442",X"0008",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"04F5",X"0442",X"0003",X"00BB",X"0164",X"06DB",X"04D0",X"0442",
X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"04CA",X"0442",X"0006",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"04E0",X"0442",X"0004",X"00BB",X"0164",
X"06DB",X"0F1B",X"01A4",X"FF00",X"0060",X"0033",X"0010",X"FFFF",
X"044C",X"000A",X"FF01",X"FF00",X"0422",X"044C",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"041E",X"044C",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"041B",X"044C",X"000A",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
X"0421",X"044C",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0060",
X"001C",X"0011",X"FFFF",X"044C",X"000A",X"FF01",X"FF00",X"0441",
X"044C",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"046F",X"044C",X"0005",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0060",X"0063",X"0012",X"FFFF",X"044C",
X"000A",X"FF01",X"FF00",X"0493",X"044C",X"000A",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
X"04A6",X"044C",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"04B2",X"044C",X"0008",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"04A2",X"044C",X"0005",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"04AD",X"044C",X"0009",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"012A",X"0499",X"044C",X"0003",X"00BB",X"0164",X"06DB",X"04AC",
X"044C",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"04BB",X"044C",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"04AB",X"044C",X"0008",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"0060",X"0048",
X"0013",X"FFFF",X"044C",X"000A",X"FF01",X"FF00",X"04D1",X"044C",
X"0003",X"00BB",X"0164",X"06DB",X"04C2",X"044C",X"0007",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"04E0",X"044C",
X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"04C7",X"044C",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"04E1",X"044C",X"0008",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"04ED",X"044C",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"04F0",X"044C",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0060",X"002E",
X"0014",X"FFFF",X"044C",X"000A",X"FF01",X"FF00",X"0429",X"044C",
X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"0417",X"044C",X"0003",X"00BB",X"0164",X"06DB",
X"0404",X"044C",X"0009",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"040A",X"044C",X"0005",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0060",X"001C",X"0015",X"FFFF",
X"044C",X"000A",X"FF01",X"FF00",X"0470",X"044C",X"0004",X"00BB",
X"0164",X"06DB",X"0F1B",X"0468",X"044C",X"000A",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
X"0060",X"0020",X"0016",X"FFFF",X"044C",X"000A",X"FF01",X"FF00",
X"04B7",X"044C",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0486",X"044C",X"0008",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",
X"0060",X"003E",X"0017",X"FFFF",X"044C",X"000A",X"FF01",X"FF00",
X"04DE",X"044C",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"04FB",X"044C",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"04F9",X"044C",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"04C7",X"044C",X"000A",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"04EC",
X"044C",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"04F3",
X"044C",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"0194",X"FF00",
X"0060",X"0049",X"0010",X"FFFF",X"0456",X"000B",X"FF01",X"FF00",
X"0403",X"0456",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0429",X"0456",X"0006",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0438",X"0456",
X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"043E",X"0456",
X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"043A",
X"0456",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"042D",X"0456",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"0435",X"0456",X"0004",X"00BB",X"0164",X"06DB",
X"0F1B",X"0060",X"002E",X"0011",X"FFFF",X"0456",X"000B",X"FF01",
X"FF00",X"0447",X"0456",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"0478",X"0456",X"000A",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0478",
X"0456",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"0459",X"0456",X"0003",X"00BB",X"0164",X"06DB",X"0060",
X"0044",X"0012",X"FFFF",X"0456",X"000B",X"FF01",X"FF00",X"0484",
X"0456",X"0003",X"00BB",X"0164",X"06DB",X"0484",X"0456",X"0007",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"0485",
X"0456",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"01E3",X"012A",X"00E0",X"04AD",X"0456",X"0006",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"04B3",X"0456",X"0006",
X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"0495",X"0456",
X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",
X"01E3",X"012A",X"00E0",X"0060",X"002E",X"0013",X"FFFF",X"0456",
X"000B",X"FF01",X"FF00",X"04CA",X"0456",X"000A",X"00BB",X"0164",
X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",X"00E0",
X"04E1",X"0456",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",X"04FD",
X"0456",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"04F8",X"0456",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"0060",X"002B",X"0014",X"FFFF",X"0456",X"000B",X"FF01",
X"FF00",X"0437",X"0456",X"0004",X"00BB",X"0164",X"06DB",X"0F1B",
X"0421",X"0456",X"0005",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"040A",X"0456",X"000A",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",
X"0607",X"036C",X"01E3",X"012A",X"00E0",X"0412",X"0456",X"0004",
X"00BB",X"0164",X"06DB",X"0F1B",X"0060",X"0008",X"0015",X"FFFF",
X"0456",X"000B",X"FF01",X"FF00",X"0060",X"004D",X"0016",X"FFFF",
X"0456",X"000B",X"FF01",X"FF00",X"048F",X"0456",X"0004",X"00BB",
X"0164",X"06DB",X"0F1B",X"04B3",X"0456",X"0003",X"00BB",X"0164",
X"06DB",X"04A2",X"0456",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"0488",X"0456",X"0003",X"00BB",X"0164",
X"06DB",X"04B6",X"0456",X"0006",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"04A1",X"0456",X"0005",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0482",X"0456",X"0007",X"00BB",X"0164",X"06DB",
X"0F1B",X"0980",X"0607",X"036C",X"04B1",X"0456",X"000A",X"00BB",
X"0164",X"06DB",X"0F1B",X"0980",X"0607",X"036C",X"01E3",X"012A",
X"00E0",X"0060",X"0029",X"0017",X"FFFF",X"0456",X"000B",X"FF01",
X"FF00",X"04FA",X"0456",X"0003",X"00BB",X"0164",X"06DB",X"04FF",
X"0456",X"0007",X"00BB",X"0164",X"06DB",X"0F1B",X"0980",X"0607",
X"036C",X"04C7",X"0456",X"0008",X"00BB",X"0164",X"06DB",X"0F1B",
X"0980",X"0607",X"036C",X"01E3",X"04E1",X"0456",X"0003",X"00BB",
X"0164",X"06DB");

Type iLinkFR_Array is Array(0 to 2) of std_logic_vector(9 downto 0);
signal iLinkFR : iLinkFR_Array;

signal LinkDCODL : std_logic_vector(1 downto 0);

signal Gap_Count : std_logic_vector(3 downto 0) := (others => '0');
signal BusTimer : std_logic_vector(4 downto 0) := (others => '0');

signal IntDCOClk,IntClk : std_logic;
signal DValid : std_logic_vector(2 downto 0);
signal IntClr : std_logic := '0';

Type CounterArray is Array(0 to 2) of std_logic_vector(15 downto 0);
signal TxCount  : CounterArray;

Type WdCntArray is Array (0 to 2) of std_logic_vector(15 downto 0);
Constant WdCnt : WdCntArray := (X"15D1",X"14E7",X"14AA");

Type Index_array is array(0 to 2) of Integer;
constant iWdCnt : Index_array := (LinkDat0_Size,LinkDat1_Size,LinkDat2_Size);

Type LinkArray is Array (0 to 71) of std_logic_vector(15 downto 0);
Constant LinkDat : LinkArray := (x"0018",x"0001",x"0021",x"0022",
                                 x"0023",x"0024",x"0025",x"0026",
											x"0027",x"0028",x"0029",x"002A",
											x"002B",x"002C",x"002D",x"002E",
											x"002F",x"0030",x"0031",x"0032",
											x"0033",x"0034",x"0035",x"0036",
											x"0018",x"0002",x"0031",x"0032",
                                 x"0033",x"0034",x"0035",x"0036",
											x"0037",x"0038",x"0039",x"003A",
                                 x"003B",x"003C",x"003D",x"003E",
											x"003F",x"0040",x"0041",x"0042",
											x"0043",x"0044",x"0045",x"0046",
											x"0018",x"0004",x"0041",x"0042",
                                 x"0043",x"0044",x"0045",x"0046",
											x"0047",x"0048",x"0049",x"004A",
                                 x"004B",x"004C",x"004D",x"004E",
											x"004F",x"0050",x"0051",x"0052",
											x"0053",x"0054",x"0055",x"0056");

Type ShiftArray is Array(0 to 2) of std_logic_vector(9 downto 0); 
signal TxReg0,TxReg1 : ShiftArray;

signal Tx1Val : std_logic_vector(15 downto 0);
signal CrCEn0,CRCRst0,CrCEn1,CRCRst1,TxWait : std_logic;
signal uCWRDL : std_logic_vector(1 downto 0);
signal MarkerCount : std_logic_vector(6 downto 0);
signal Clk53Mhz,Marker,Even_Odd,MarkerReq,Clk160Mhz : std_logic;
signal BunchBits : std_logic_vector(3 downto 0); 
signal BunchCount : std_logic_vector(2 downto 0); 

-- signal PeriodicMicrobunch, IntTmgEn: std_logic;

begin

-- Instantiate the Unit Under Test (UUT)
uut: ControllerFPGA_1 
	PORT MAP 
	(VXO_P => VXO_P,VXO_N => VXO_N,ClkB_P => ClkB_P,ClkB_N => ClkB_N,
	 Clk50MHz => Clk50MHz,BnchClk => BnchClk,
-- 156.25 MHz GTP Reference clock, Gigabit data lines
	GTPClk_P => GTPClk_P,GTPClk_N => GTPClk_N,GTPRx_P => GTPRx_P,
	GTPRx_N => GTPRx_N, GTPTx_P => GTPTx_P, GTPTx_N => GTPTx_N,
	TDisA => TDisA,TDisB => TDisB,
	SD_A => SD_A,SD_B => SD_B,
	CpldRst => CpldRst, CpldCS => CpldCS, uCRd => uCRd, 
	uCWr => uCWr, EthCS => EthCS,
	uCA => uCA,	uCD => uCD, GA => GA,
	LINKClk_P => LINKClk_P,LINKClk_N => LINKClk_N,
	LinkFR_P => LinkFR_P,LinkFR_N => LinkFR_N,
	LinkSDat_P => LinkSDat_P,LinkSDat_N => LinkSDat_N,
	HeartBeatFM => HeartBeatFM,TrigFM => TrigFM,
	uBunchLED => uBunchLED,TrigLED => TrigLED,
	PllSClk => PllSClk,PllSDat => PllSDat,PllLd => PllLd,
	PllPDn => PllPDn, PllStat => PllStat,
	LEDSClk => LEDSClk,LEDSDat => LEDSDat,
	LEDLd => LEDLd, LEDRst => LEDRst,
	DQ => DQ, ZEthA => ZEthA, ZEthCS => ZEthCS,
	ZEthWE => ZEthWE,ZEthClk => ZEthClk,
	ZEthBE => ZEthBE,	ZEthEOF => ZEthEOF,
	ZEthLen => ZEthLen, GPO => GPO,
	GPI => GPI,NimTrig => NimTrig,
	-- PeriodicMicrobunch => PeriodicMicrobunch, IntTmgEn => IntTmgEn,
	Debug => Debug);

--TxCRCGEn : crc 
-- port map( data_in => uCD,
--    crc_en => CrCEn0, rst => CRCRst0, clk => GTPClk_P(0),
--    crc_out => TxCRC0);
--
--CRCRst0 <= '1' when uCA <= "00" & GTPWrtAddr(0) and uCWR = '0' and CpldCS = '0' else '0';
--
--CRCRst1 <= '1' when uCA <= "00" & GTPWrtAddr(2) and uCWR = '0' and CpldCS = '0' else '0';

-- Cross connect GTP I/O for loopback operation
-- Rx0 input polarity is inverted
--GTPRx_N(0) <= GTPTx_P(1);
--GTPRx_P(0) <= GTPTx_N(1);

GTPRx_N(1) <= GTPTx_N(0);
GTPRx_P(1) <= GTPTx_P(0);

Init_Process : process
	begin
		CpldRst <= '0'; GA <= "00";
		TxWait <= '0';
		wait for 100 ns;
		CpldRst <= '1';
		wait for 1 us;
		TxWait <= '1';
	wait;
	end process;

-- Clock process definitions

-- Generate a 1695 ns interval
Clk53Mhz_Process : process
   begin
		Clk53Mhz <= '0'; 
		wait for Clk53Mhz_Period/2;
		Clk53Mhz <= '1'; 
		wait for Clk53Mhz_Period/2;
   end process;

-- Encoded Bunch clock
Clk160Mhz_Process : process
   begin
		Clk160Mhz <= '0'; 
		wait for Clk160Mhz_Period/2;
		Clk160Mhz <= '1'; 
		wait for Clk160Mhz_Period/2;
   end process;

-- 100 Mhz System Clocks
ClkB_P_process :process
   begin
		ClkB_P <= '0'; VXO_P <= '0'; 
		ClkB_N <= '1'; VXO_N <= '1'; 
		wait for ClkB_P_period/2;
		ClkB_P <= '1'; VXO_P <= '1'; 
		ClkB_N <= '0'; VXO_N <= '0'; 
		wait for ClkB_P_period/2;
   end process;

Clk50MhzProcess : process
    begin
	  Clk50MHz <= '0';
	  wait for Clk50Mhz_Period/2;
	  Clk50MHz <= '1';
	  wait for Clk50Mhz_Period/2;
	 end process;

GTP_Ref_Clk_process :process
   begin
		GTPClk_P <= "00"; GTPClk_N <= "11"; 
		wait for GTPRefClk_Period/2;
		GTPClk_P <= "11"; GTPClk_N <= "00"; 
		wait for GTPRefClk_Period/2;
   end process;

LINK_Clk_process : process
  begin
	LINKClk_P <= "000";
	LINKClk_N <= "111";
	 wait for DCO_period/2;
	LINKClk_P <= "111";
	LINKClk_N <= "000";
	 wait for DCO_period/2;
   end process;

IntClk_Clk_process : process
  begin
	IntClk <= '0';
	 wait for DCO_period * 2.5;
	IntClk <= '1';
	 wait for DCO_period * 2.5;
   end process;

-- Generate a marker every 90 RF ticks
Marker_Process : process(CpldRst,Clk53Mhz)

begin

	if CpldRst = '0' then
		
		MarkerCount <= (others => '0');
		Marker <= '0'; Even_Odd <= '0';

	elsif rising_edge (Clk53Mhz) then

		  if MarkerCount /= 89 then MarkerCount <= MarkerCount + 1;
		  else MarkerCount <= (others => '0');
		  end if;

		  if MarkerCount = 89 then 
				Marker <= '1';
				Even_Odd <= not Even_Odd;
		  elsif MarkerReq = '1' 
				then Marker <= '0';
				Even_Odd <= Even_Odd;
		  else
				Marker <= Marker;
				Even_Odd <= Even_Odd;
		  end if;

   end if; -- CpldRst;

end process;

Bunch_process : process(CpldRst,Clk160Mhz)

 begin

  if CpldRst = '0' then

	 BunchBits <= X"C"; BunchCount <= "000";
	 MarkerReq <= '0';

   elsif rising_edge(Clk160Mhz) then

		if ((MarkerReq = '0' and BunchCount = 3)
		 or (MarkerReq = '1' and BunchCount = 7)) then BunchCount <= "000";
		else BunchCount <= BunchCount + 1;
		end if;

		if MarkerReq = '0' and Marker = '1' and BunchCount = 3 then MarkerReq <= '1';
		 elsif MarkerReq = '1' and BunchCount = X"7"
		   then MarkerReq <= '0';
		 else MarkerReq <= MarkerReq;
		end if;

		Case Even_Odd is 
		 when '0' =>
			   if (MarkerReq = '0' and (BunchCount = 0 or BunchCount = 1))
				or (MarkerReq = '1' and (BunchCount = 0 or BunchCount = 4 or BunchCount = 5 or BunchCount = 6))
			  then BnchClk <= '1'; 
			else BnchClk <= '0';
			end if;
		 when '1' =>
			   if (MarkerReq = '0' and (BunchCount = 0 or BunchCount = 1))
				or (MarkerReq = '1' and (BunchCount = 0 or BunchCount = 1 or BunchCount = 2 or BunchCount = 4))
			  then BnchClk <= '1'; 
			else BnchClk <= '0';
			end if;
		  when others => BnchClk <= '0'; 
		 end case;
		 
 end if; -- CpldRst

end process;

-- Stimulus process

-- Clk0    -_-_-_-_-_-_-_-_-_-_
-- Frame0  -----_____-----_____
-- Lane 01 V1DDDV1dddV1DDDV1ddd
-- Lane 00 DDDDDdddddDDDDDddddd

-- Clk1    -_-_-_-_-_-_-_-_-_-_
-- Frame1  _____-----_____-----
-- Lane 11 V1DDDV1dddV1DDDV1ddd
-- Lane 10 DDDDDdddddDDDDDddddd

-- Clk2    -_-_-_-_-_-_-_-_-_-_
-- Frame2  -----_____-----_____
-- Lane 21 V1DDDV1dddV1DDDV1ddd
-- Lane 20 DDDDDdddddDDDDDddddd

shift_proc: process(CpldRst,LINKClk_P(0))

Variable Index : Index_array;

begin

if CpldRst = '0' then
	LinkDCODL <= "00";
	iLinkFR <= (others => ("00" & X"1F"));
	LinkSDat_P <= (others => '0');
	LinkSDat_N <= (others => '1');
	DValid <= "000";
	Index(0) := 0; Index(1) := 0; Index(2) := 0;
	TxReg1 <= (others => (others => '0'));
	TxReg0 <= (others => (others => '0'));
	TxCount <= (others => X"0000");

elsif (LINKClk_P(0)' event)

  then

	LinkDCODL(0) <= IntClk;
	LinkDCODL(1) <= LinkDCODL(0);
	
for i in 0 to 2 loop

	if LinkDCODL = "01" then 
	if DValid(i) = '1' and TxCount(i) /= WdCnt(i) then TxCount(i) <= TxCount(i) + 1;
	elsif DValid(i) = '1' and TxCount(i) = WdCnt(i) then TxCount(i) <= X"0000";
	else TxCount(i) <= TxCount(i);
	end if;
	end if;

end loop;

	if LinkDCODL = "01" and Index(0) < iWdCnt(0) then 
-- The framing signal is high at the beginning of the serial word
    iLinkFR(0) <= "11" & X"E0";
-- Locad a data value
	 TxReg1(0) <= DValid(0) & '1' & LinkDat0(Index(0))(15 downto 13) & DValid(0) & '1' & LinkDat0(Index(0))(7 downto 5);
	 TxReg0(0) <= LinkDat0(Index(0))(12 downto 8) & LinkDat0(Index(0))(4 downto 0);
--  then shift out
	else 
	 TxReg1(0) <= TxReg1(0)(8 downto 0) & '0';
	 TxReg0(0) <= TxReg0(0)(8 downto 0) & '0';
	 iLinkFR(0) <= iLinkFR(0)(8 downto 0) & iLinkFR(0)(9);
	end if;

	if LinkDCODL = "01" and Index(1) < iWdCnt(1) then 
-- The framing signal is high at the beginning of the serial word
    iLinkFR(1) <= "11" & X"E0";
-- Locad a data value
	 TxReg1(1) <= DValid(1) & '1' & LinkDat1(Index(1))(15 downto 13) & DValid(1) & '1' & LinkDat1(Index(1))(7 downto 5);
	 TxReg0(1) <= LinkDat1(Index(1))(12 downto 8) & LinkDat1(Index(1))(4 downto 0);
--  then shift out
	else 
	 TxReg1(1) <= TxReg1(1)(8 downto 0) & '0';
	 TxReg0(1) <= TxReg0(1)(8 downto 0) & '0';
	 iLinkFR(1) <= iLinkFR(1)(8 downto 0) & iLinkFR(1)(9);
	end if;

	if LinkDCODL = "01" and Index(2) < iWdCnt(2) then 
-- The framing signal is high at the beginning of the serial word
    iLinkFR(2) <=  "11" & X"E0";
-- Locad a data value
	 TxReg1(2) <= DValid(2) & '1' & LinkDat2(Index(2))(15 downto 13) & DValid(2) & '1' & LinkDat2(Index(2))(7 downto 5);
	 TxReg0(2) <= LinkDat2(Index(2))(12 downto 8) & LinkDat2(Index(2))(4 downto 0);
--  then shift out
	else 
	 TxReg1(2) <= TxReg1(2)(8 downto 0) & '0';
	 TxReg0(2) <= TxReg0(2)(8 downto 0) & '0';
	 iLinkFR(2) <= iLinkFR(2)(8 downto 0) & iLinkFR(2)(9);
	end if;

for i in 0 to 2 loop

	if LinkDCODL = "10" and DValid(i) = '1' and Index(i) /= iWdCnt(i)
		then Index(i) := Index(i) + 1;
	else Index(i) := Index(i); 
	end if;

if i = 0
then
	if TxWait = '1' and DValid(i) <= '0' and TxCount(i) /= WdCnt(i) then DValid(i) <= '1';
	 elsif LinkDCODL = "10" and DValid(i) <= '1' and TxCount(i) = WdCnt(i) then DValid(i) <= '0';
	 else DValid(i) <= DValid(i);
	end if;
else
	 DValid(i) <= '0';
end if;

LinkSDat_P(2*i+1) <=     TxReg1(i)(9) after 0.5 ns;
LinkSDat_N(2*i+1) <= not TxReg1(i)(9) after 0.5 ns;

LinkSDat_P(2*i) <=     TxReg0(i)(9) after 0.5 ns;
LinkSDat_N(2*i) <= not TxReg0(i)(9) after 0.5 ns;

if i = 1
then
LinkFR_N(i) <=     iLinkFR(i)(9) after 0.5 ns;
LinkFR_P(i) <= not iLinkFR(i)(9) after 0.5 ns;
else
LinkFR_P(i) <=     iLinkFR(i)(9) after 0.5 ns;
LinkFR_N(i) <= not iLinkFR(i)(9) after 0.5 ns;

end if;

end loop;

end if;

end process;


-- DG: external trigger process
Trigger: process
begin
NimTrig <= '0';

wait for 4000 ns;
-- send a trigger -- OFF beam
NimTrig <= '1';
wait for 25 ns;
NimTrig <= '0';

wait;-- for 300 ns;

--
---- send a trigger -- ON beam
--NimTrig <= '1';
--wait for 200 ns;
--NimTrig <= '0';
--
--wait for 300 ns;
--
---- send a trigger -- ON beam
--NimTrig <= '1';
--wait for 200 ns;
--NimTrig <= '0';

end process;

-- DG: PPS process
PPS: process
begin
GPI <= '0';
wait for 1 us;
GPI <= '1';
wait for 100 ns;
GPI <= '0';
end process;


uCIO : process

		Variable GIndex : integer range 0 to GTP_Size - 1;

	begin
		uCWr <= '1'; uCRd <= '1';
		uCA <= (Others => 'Z');
		uCD <= (others => 'Z'); 
		CpldCS <= '1'; EthCS <= '1';
		Tx1Val <= X"1111";

	wait for 1 us;	

		  uCA <= "00" & ActvRegAddrHi;
		  wait for 5 ns;
		  CpldCS <= '0';
		  wait for 5 ns;
		  uCD <= X"0000";
		  uCWr <= '0';
		  wait for 15 ns;
		  uCWr <= '1';
		  CpldCS <= '1';
		  wait for 5 ns;
		  uCA <= (Others => 'Z');
		  uCD <= (others => 'Z');
		  wait for 10 ns;
	wait for 100 ns;	

		  uCA <= "00" & ActvRegAddrLo;
		  wait for 5 ns;
		  CpldCS <= '0';
		  wait for 5 ns;
		  uCD <= X"0101";
		  uCWr <= '0';
		  wait for 15 ns;
		  uCWr <= '1';
		  CpldCS <= '1';
		  wait for 5 ns;
		  uCA <= (Others => 'Z');
		  uCD <= (others => 'Z');
		  wait for 10 ns;
	wait for 100 ns;	

		  uCA <= "00" & DReqBrstCntAd;
		  wait for 5 ns;
		  CpldCS <= '0';
		  wait for 5 ns;
		  uCD <= X"0005";
		  uCWr <= '0';
		  wait for 15 ns;
		  uCWr <= '1';
		  CpldCS <= '1';
		  wait for 5 ns;
		  uCA <= (Others => 'Z');
		  uCD <= (others => 'Z');
		  wait for 10 ns;

	wait for 100 ns;	

		  uCA <= "00" & HrtBtBrstCntAdLo;
		  wait for 5 ns;
		  CpldCS <= '0';
		  wait for 5 ns;
		  uCD <= X"0100";
		  uCWr <= '0';
		  wait for 15 ns;
		  uCWr <= '1';
		  CpldCS <= '1';
		  wait for 5 ns;
		  uCA <= (Others => 'Z');
		  uCD <= (others => 'Z');
		  wait for 10 ns;

	wait for 1 us;	

		  uCA <= "00" & CSRRegAddr;
		  wait for 5 ns;
		  CpldCS <= '0';
		  wait for 5 ns;
--		  uCD <= X"0040";
			-- turns on IntTmgEn and TstTrigEn
		  uCD <= X"0101";
--		  uCD <= X"0303";
		  uCWr <= '0';
		  wait for 15 ns;
		  uCWr <= '1';
		  CpldCS <= '1';
		  wait for 5 ns;
		  uCA <= (Others => 'Z');
		  uCD <= (others => 'Z');
		  wait for 10 ns;
		  
	wait for 200 ns;
		  uCA <= "00" & ExternalTriggerControlAddress;
		  wait for 5 ns;
		  CpldCS <= '0';
		  wait for 5 ns;
		  -- Periodic Microbunch ON, reset Ext Trig timestamp ON, Pulse detect gate 15	
		  uCD <= X"00FC";
		  uCWr <= '0';
		  wait for 15 ns;
		  uCWr <= '1';
		  CpldCS <= '1';
		  wait for 5 ns;
		  uCA <= (Others => 'Z');
		  uCD <= (others => 'Z');
		  wait for 10 ns;	
	wait for 50 ns;
		  uCA <= "00" & PeriodicMicrobunchPeriodAddrLo;
		  wait for 5 ns;
		  CpldCS <= '0';
		  wait for 5 ns;
		  uCD <= X"000F";
		  uCWr <= '0';
		  wait for 15 ns;
		  uCWr <= '1';
		  CpldCS <= '1';
		  wait for 5 ns;
		  uCA <= (Others => 'Z');
		  uCD <= (others => 'Z');
		  wait for 10 ns;	
		  
	-- turn external trigger generation of microbunches back on
	wait for 500 ns;
		  uCA <= "00" & ExternalTriggerControlAddress;
		  wait for 5 ns;
		  CpldCS <= '0';
		  wait for 5 ns;
		  -- Periodic Microbunch OFF, reset Ext Trig timestamp ON, Pulse detect gate 15	
		  uCD <= X"00F8";
		  uCWr <= '0';
		  wait for 15 ns;
		  uCWr <= '1';
		  CpldCS <= '1';
		  wait for 5 ns;
		  uCA <= (Others => 'Z');
		  uCD <= (others => 'Z');
		  wait for 10 ns;	
	-- start inhibit triggers
	wait for 100 ns;
		uCA <= "00" & ExternalTriggerInhibitAddrLo;
		  wait for 5 ns;
		  CpldCS <= '0';
		  wait for 5 ns;
		  uCD <= X"003C";
		  uCWr <= '0';
		  wait for 15 ns;
		  uCWr <= '1';
		  CpldCS <= '1';
		  wait for 5 ns;
		  uCA <= (Others => 'Z');
		  uCD <= (others => 'Z');
		  wait for 10 ns;	
		  
	wait for 100 ns;
			uCA <= "00" & PLLHiAddr;
		  wait for 5 ns;
		  CpldCS <= '0';
		  wait for 5 ns;
		  uCD <= X"0000";
		  uCWr <= '0';
		  wait for 25 ns;
		  uCWr <= '1';
		  CpldCS <= '1';
		  wait for 5 ns;
		  uCA <= (Others => 'Z');
		  uCD <= (others => 'Z');
		  wait for 10 ns;	
		  
	wait for 50 ns;
		  		uCA <= "00" & PLLLoAddr;
		  wait for 5 ns;
		  CpldCS <= '0';
		  wait for 5 ns;
		  uCD <= X"0008";
		  uCWr <= '0';
		  wait for 25 ns;
		  uCWr <= '1';
		  CpldCS <= '1';
		  wait for 5 ns;
		  uCA <= (Others => 'Z');
		  uCD <= (others => 'Z');
		  wait for 10 ns;	
		  
	wait for 50 ns;

		  		uCA <= "00" & PLLLoAddr;
		  wait for 5 ns;
		  CpldCS <= '0';
		  wait for 5 ns;
		  uCD <= X"0051";
		  uCWr <= '0';
		  wait for 25 ns;
		  uCWr <= '1';
		  CpldCS <= '1';
		  wait for 5 ns;
		  uCA <= (Others => 'Z');
		  uCD <= (others => 'Z');
		  wait for 10 ns;	
		  
  wait for 2500 ns;
		uCA <= "00" & TRigReqBuffAd;
		  uCD <= (others => 'Z');

		  wait for 5 ns;
		  CpldCS <= '0';
		  wait for 10 ns;
		  uCRD <= '0';
		  wait for 50 ns;
		  uCRD <= '1';
		  CpldCS <= '1';
		  wait for 10 ns;
		  uCA <= (Others => 'Z');
		  wait for 50 ns;
			

		  uCA <= "00" & TRigReqBuffAd;
		  wait for 5 ns;
		  CpldCS <= '0';
		  wait for 10 ns;
		  uCRD <= '0';
		  wait for 50 ns;
		  uCRD <= '1';
		  CpldCS <= '1';
		  wait for 10 ns;
		  uCA <= (Others => 'Z');
		  wait for 50 ns;
		  		uCA <= "00" & TRigReqBuffAd;
		  wait for 5 ns;
		  CpldCS <= '0';
		  wait for 10 ns;
		  uCRD <= '0';
		  wait for 50 ns;
		  uCRD <= '1';
		  CpldCS <= '1';
		  wait for 10 ns;
		  uCA <= (Others => 'Z');
		  wait for 50 ns;
		
--
--	wait for 1 us;	

-- Send the packet preamble

--		  uCA <= "00" & GTPWrtAddr(1);
-- 		  wait for 5 ns;
--		  CpldCS <= '0';
--		  wait for 5 ns;
--		  uCD <= X"0002";
--		  uCWr <= '0';
--		  wait for 15 ns;
--		  uCWr <= '1';
--		  CpldCS <= '1';
--		  wait for 5 ns;
--		  uCA <= (Others => 'Z');
--		  uCD <= (others => 'Z');
--		  wait for 10 ns;

--		  uCA <= "00" & GTPWrtAddr(0);
-- 	  wait for 5 ns;
--		  CpldCS <= '0';
--		  wait for 5 ns;
--		  uCD <= X"0003";
--		  uCWr <= '0';
--		  wait for 15 ns;
--		  uCWr <= '1';
--		  EthCS <= '1';
--		  wait for 5 ns;
--		  uCA <= (Others => 'Z');
--		  uCD <= (others => 'Z');
--		  wait for 10 ns;

--for GIndex in 0 to 7 loop
 
-- Send the packet body
--		  uCA <= "00" & GTPWrtAddr(3);
-- 		  wait for 5 ns;
--		  CpldCS <= '0';
--		  wait for 5 ns;
--		  uCD <= TxVal(GIndex);
--		  uCWr <= '0';
--		  wait for 15 ns;
--		  uCWr <= '1';
--		  CpldCS <= '1';
--		  wait for 5 ns;
--		  uCA <= (Others => 'Z');
--		  uCD <= (others => 'Z');
--		  wait for 10 ns;

--		  uCA <= "00" & GTPWrtAddr(2);
-- 	  wait for 5 ns;
--		  CpldCS <= '0';
--		  wait for 5 ns;
--		  uCD <= Tx1Val;
--		  uCWr <= '0';
--		  wait for 15 ns;
--		  uCWr <= '1';
--		  EthCS <= '1';
--		  wait for 5 ns;
--		  uCA <= (Others => 'Z');
--		  uCD <= (others => 'Z');
--		  wait for 10 ns;

--		  Tx1Val <= Tx1Val + X"1111";

--		end loop;

-- Send the packet CRC

--		  uCA <= "00" & GTPWrtAddr(5);
-- 		  wait for 5 ns;
--		  CpldCS <= '0';
--		  wait for 5 ns;
--		  uCD <= X"0002";
--		  uCWr <= '0';
--		  wait for 15 ns;
--		  uCWr <= '1';
--		  CpldCS <= '1';
--		  wait for 5 ns;
--		  uCA <= (Others => 'Z');
--		  uCD <= (others => 'Z');
--		  wait for 10 ns;

--		  uCA <= "00" & GTPWrtAddr(5);
-- 	  wait for 5 ns;
--		  CpldCS <= '0';
--		  wait for 5 ns;
--		  uCD <= X"0003";
--		  uCWr <= '0';
--		  wait for 15 ns;
--		  uCWr <= '1';
--		  EthCS <= '1';
--		  wait for 5 ns;
--		  uCA <= (Others => 'Z');
--		  uCD <= (others => 'Z');
--		  wait for 10 ns;
	
--		  uCA <= "00" & GTPRdAddr0;
-- 		  wait for 5 ns;
--		  CpldCS <= '0';
--		  wait for 10 ns;
--		  uCRD <= '0';
--		  wait for 50 ns;
--		  uCRD <= '1';
--		  CpldCS <= '1';
--		  wait for 10 ns;
--		  uCA <= (Others => 'Z');
--		  wait for 50 ns;

--		  uCA <= "00" & GTPRdAddr1;
-- 		  wait for 5 ns;
--		  CpldCS <= '0';
--		  wait for 10 ns;
--		  uCRD <= '0';
--		  wait for 30 ns;
--		  uCRD <= '1';
--		  CpldCS <= '1';
--		  wait for 10 ns;
--		  uCA <= (Others => 'Z');
--		  wait for 50 ns;

		  wait;

end process uCIO;

DQIO : process


	begin
		DQ <= (others => 'Z'); 
		
	wait for 2859 ns;	

	DQ <= X"1234";  
	
	wait for 15 ns;
	
		DQ <= (others => 'Z'); 
	wait;

end process DQIO;

END;
